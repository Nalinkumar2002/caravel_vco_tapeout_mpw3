magic
tech sky130A
magscale 1 2
timestamp 1635398265
<< nwell >>
rect -36844 43530 -35986 45134
rect -36846 42976 -35986 43530
rect -36850 42720 -35986 42976
rect -36850 42592 -35988 42720
<< nmos >>
rect -37134 44878 -37004 44914
rect -37292 44600 -37004 44636
rect -37582 44184 -37324 44220
rect -37106 44184 -37006 44220
rect -37582 43912 -37324 43948
rect -37106 43912 -37006 43948
rect -37582 43640 -37324 43676
rect -37106 43640 -37006 43676
rect -37582 43368 -37324 43404
rect -37108 43368 -37008 43404
rect -37582 43096 -37324 43132
rect -37108 43096 -37008 43132
rect -37524 42766 -37322 42802
<< pmos >>
rect -36790 44878 -36532 44914
rect -36790 44600 -36214 44636
rect -36790 44184 -36690 44220
rect -36478 44186 -36218 44222
rect -36790 43912 -36690 43948
rect -36478 43914 -36218 43950
rect -36790 43640 -36690 43676
rect -36478 43642 -36218 43678
rect -36792 43368 -36692 43404
rect -36478 43370 -36218 43406
rect -36792 43096 -36692 43132
rect -36478 43098 -36218 43134
rect -36478 42764 -36276 42800
<< ndiff >>
rect -37134 44986 -37004 45004
rect -37134 44950 -37074 44986
rect -37038 44950 -37004 44986
rect -37134 44914 -37004 44950
rect -37134 44842 -37004 44878
rect -37134 44806 -37074 44842
rect -37038 44806 -37004 44842
rect -37134 44788 -37004 44806
rect -37292 44708 -37004 44726
rect -37292 44672 -37268 44708
rect -37234 44672 -37194 44708
rect -37160 44672 -37126 44708
rect -37092 44672 -37056 44708
rect -37020 44672 -37004 44708
rect -37292 44636 -37004 44672
rect -37292 44564 -37004 44600
rect -37292 44528 -37268 44564
rect -37234 44528 -37194 44564
rect -37160 44528 -37126 44564
rect -37092 44528 -37058 44564
rect -37022 44528 -37004 44564
rect -37292 44510 -37004 44528
rect -37582 44292 -37324 44310
rect -37582 44256 -37552 44292
rect -37518 44256 -37478 44292
rect -37444 44256 -37398 44292
rect -37364 44256 -37324 44292
rect -37106 44292 -37006 44310
rect -37106 44256 -37074 44292
rect -37038 44256 -37006 44292
rect -37582 44220 -37324 44256
rect -37106 44220 -37006 44256
rect -37582 44150 -37324 44184
rect -37582 44148 -37398 44150
rect -37582 44112 -37552 44148
rect -37516 44112 -37476 44148
rect -37440 44114 -37398 44148
rect -37364 44114 -37324 44150
rect -37440 44112 -37324 44114
rect -37582 44094 -37324 44112
rect -37106 44148 -37006 44184
rect -37106 44112 -37074 44148
rect -37038 44112 -37006 44148
rect -37106 44094 -37006 44112
rect -37582 44020 -37324 44038
rect -37582 43984 -37552 44020
rect -37518 43984 -37478 44020
rect -37444 43984 -37398 44020
rect -37364 43984 -37324 44020
rect -37106 44020 -37006 44038
rect -37106 43984 -37074 44020
rect -37038 43984 -37006 44020
rect -37582 43948 -37324 43984
rect -37106 43948 -37006 43984
rect -37582 43878 -37324 43912
rect -37582 43876 -37398 43878
rect -37582 43840 -37552 43876
rect -37516 43840 -37476 43876
rect -37440 43842 -37398 43876
rect -37364 43842 -37324 43878
rect -37440 43840 -37324 43842
rect -37582 43822 -37324 43840
rect -37106 43876 -37006 43912
rect -37106 43840 -37074 43876
rect -37038 43840 -37006 43876
rect -37106 43822 -37006 43840
rect -37582 43748 -37324 43766
rect -37582 43712 -37552 43748
rect -37518 43712 -37478 43748
rect -37444 43712 -37398 43748
rect -37364 43712 -37324 43748
rect -37106 43748 -37006 43766
rect -37106 43712 -37074 43748
rect -37038 43712 -37006 43748
rect -37582 43676 -37324 43712
rect -37106 43676 -37006 43712
rect -37582 43606 -37324 43640
rect -37582 43604 -37398 43606
rect -37582 43568 -37552 43604
rect -37516 43568 -37476 43604
rect -37440 43570 -37398 43604
rect -37364 43570 -37324 43606
rect -37440 43568 -37324 43570
rect -37582 43550 -37324 43568
rect -37106 43604 -37006 43640
rect -37106 43568 -37074 43604
rect -37038 43568 -37006 43604
rect -37106 43550 -37006 43568
rect -37582 43476 -37324 43494
rect -37582 43440 -37552 43476
rect -37518 43440 -37478 43476
rect -37444 43440 -37398 43476
rect -37364 43440 -37324 43476
rect -37108 43476 -37008 43494
rect -37108 43440 -37076 43476
rect -37040 43440 -37008 43476
rect -37582 43404 -37324 43440
rect -37108 43404 -37008 43440
rect -37582 43334 -37324 43368
rect -37582 43332 -37398 43334
rect -37582 43296 -37552 43332
rect -37516 43296 -37476 43332
rect -37440 43298 -37398 43332
rect -37364 43298 -37324 43334
rect -37440 43296 -37324 43298
rect -37582 43278 -37324 43296
rect -37108 43332 -37008 43368
rect -37108 43296 -37076 43332
rect -37040 43296 -37008 43332
rect -37108 43278 -37008 43296
rect -37582 43204 -37324 43222
rect -37582 43168 -37552 43204
rect -37518 43168 -37478 43204
rect -37444 43168 -37398 43204
rect -37364 43168 -37324 43204
rect -37108 43204 -37008 43222
rect -37108 43168 -37076 43204
rect -37040 43168 -37008 43204
rect -37582 43132 -37324 43168
rect -37108 43132 -37008 43168
rect -37582 43062 -37324 43096
rect -37582 43060 -37398 43062
rect -37582 43024 -37552 43060
rect -37516 43024 -37476 43060
rect -37440 43026 -37398 43060
rect -37364 43026 -37324 43062
rect -37440 43024 -37324 43026
rect -37582 43006 -37324 43024
rect -37108 43060 -37008 43096
rect -37108 43024 -37076 43060
rect -37040 43024 -37008 43060
rect -37108 43006 -37008 43024
rect -37524 42874 -37322 42892
rect -37524 42838 -37482 42874
rect -37448 42838 -37398 42874
rect -37364 42838 -37322 42874
rect -37524 42802 -37322 42838
rect -37524 42730 -37322 42766
rect -37524 42694 -37480 42730
rect -37444 42694 -37398 42730
rect -37362 42694 -37322 42730
rect -37524 42676 -37322 42694
<< pdiff >>
rect -36790 44986 -36532 45004
rect -36790 44950 -36758 44986
rect -36722 44950 -36686 44986
rect -36650 44950 -36616 44986
rect -36580 44950 -36532 44986
rect -36790 44914 -36532 44950
rect -36790 44842 -36532 44878
rect -36790 44806 -36758 44842
rect -36722 44806 -36688 44842
rect -36652 44806 -36618 44842
rect -36582 44806 -36532 44842
rect -36790 44788 -36532 44806
rect -36790 44710 -36214 44726
rect -36790 44708 -36688 44710
rect -36790 44672 -36758 44708
rect -36722 44674 -36688 44708
rect -36652 44674 -36618 44710
rect -36582 44674 -36548 44710
rect -36512 44674 -36478 44710
rect -36442 44674 -36408 44710
rect -36372 44674 -36338 44710
rect -36302 44674 -36268 44710
rect -36232 44674 -36214 44710
rect -36722 44672 -36214 44674
rect -36790 44636 -36214 44672
rect -36790 44564 -36214 44600
rect -36790 44528 -36758 44564
rect -36722 44528 -36688 44564
rect -36652 44528 -36618 44564
rect -36582 44528 -36548 44564
rect -36512 44528 -36478 44564
rect -36442 44528 -36408 44564
rect -36372 44528 -36338 44564
rect -36302 44528 -36268 44564
rect -36232 44528 -36214 44564
rect -36790 44510 -36214 44528
rect -36790 44292 -36690 44310
rect -36790 44256 -36758 44292
rect -36722 44256 -36690 44292
rect -36478 44294 -36218 44312
rect -36478 44258 -36436 44294
rect -36402 44258 -36356 44294
rect -36322 44258 -36282 44294
rect -36248 44258 -36218 44294
rect -36790 44220 -36690 44256
rect -36478 44222 -36218 44258
rect -36790 44148 -36690 44184
rect -36790 44112 -36758 44148
rect -36722 44112 -36690 44148
rect -36790 44094 -36690 44112
rect -36478 44152 -36218 44186
rect -36478 44116 -36436 44152
rect -36402 44150 -36218 44152
rect -36402 44116 -36360 44150
rect -36478 44114 -36360 44116
rect -36324 44114 -36284 44150
rect -36248 44114 -36218 44150
rect -36478 44096 -36218 44114
rect -36790 44020 -36690 44038
rect -36790 43984 -36758 44020
rect -36722 43984 -36690 44020
rect -36478 44022 -36218 44040
rect -36478 43986 -36436 44022
rect -36402 43986 -36356 44022
rect -36322 43986 -36282 44022
rect -36248 43986 -36218 44022
rect -36790 43948 -36690 43984
rect -36478 43950 -36218 43986
rect -36790 43876 -36690 43912
rect -36790 43840 -36758 43876
rect -36722 43840 -36690 43876
rect -36790 43822 -36690 43840
rect -36478 43880 -36218 43914
rect -36478 43844 -36436 43880
rect -36402 43878 -36218 43880
rect -36402 43844 -36360 43878
rect -36478 43842 -36360 43844
rect -36324 43842 -36284 43878
rect -36248 43842 -36218 43878
rect -36478 43824 -36218 43842
rect -36790 43748 -36690 43766
rect -36790 43712 -36758 43748
rect -36722 43712 -36690 43748
rect -36478 43750 -36218 43768
rect -36478 43714 -36436 43750
rect -36402 43714 -36356 43750
rect -36322 43714 -36282 43750
rect -36248 43714 -36218 43750
rect -36790 43676 -36690 43712
rect -36478 43678 -36218 43714
rect -36790 43604 -36690 43640
rect -36790 43568 -36758 43604
rect -36722 43568 -36690 43604
rect -36790 43550 -36690 43568
rect -36478 43608 -36218 43642
rect -36478 43572 -36436 43608
rect -36402 43606 -36218 43608
rect -36402 43572 -36360 43606
rect -36478 43570 -36360 43572
rect -36324 43570 -36284 43606
rect -36248 43570 -36218 43606
rect -36478 43552 -36218 43570
rect -36792 43476 -36692 43494
rect -36792 43440 -36760 43476
rect -36724 43440 -36692 43476
rect -36478 43478 -36218 43496
rect -36478 43442 -36436 43478
rect -36402 43442 -36356 43478
rect -36322 43442 -36282 43478
rect -36248 43442 -36218 43478
rect -36792 43404 -36692 43440
rect -36478 43406 -36218 43442
rect -36792 43332 -36692 43368
rect -36792 43296 -36760 43332
rect -36724 43296 -36692 43332
rect -36792 43278 -36692 43296
rect -36478 43336 -36218 43370
rect -36478 43300 -36436 43336
rect -36402 43334 -36218 43336
rect -36402 43300 -36360 43334
rect -36478 43298 -36360 43300
rect -36324 43298 -36284 43334
rect -36248 43298 -36218 43334
rect -36478 43280 -36218 43298
rect -36792 43204 -36692 43222
rect -36792 43168 -36760 43204
rect -36724 43168 -36692 43204
rect -36478 43206 -36218 43224
rect -36478 43170 -36436 43206
rect -36402 43170 -36356 43206
rect -36322 43170 -36282 43206
rect -36248 43170 -36218 43206
rect -36792 43132 -36692 43168
rect -36478 43134 -36218 43170
rect -36792 43060 -36692 43096
rect -36792 43024 -36760 43060
rect -36724 43024 -36692 43060
rect -36792 43006 -36692 43024
rect -36478 43064 -36218 43098
rect -36478 43028 -36436 43064
rect -36402 43062 -36218 43064
rect -36402 43028 -36360 43062
rect -36478 43026 -36360 43028
rect -36324 43026 -36284 43062
rect -36248 43026 -36218 43062
rect -36478 43008 -36218 43026
rect -36478 42874 -36276 42890
rect -36478 42872 -36376 42874
rect -36478 42836 -36446 42872
rect -36410 42838 -36376 42872
rect -36340 42838 -36276 42874
rect -36410 42836 -36276 42838
rect -36478 42800 -36276 42836
rect -36478 42728 -36276 42764
rect -36478 42692 -36436 42728
rect -36400 42692 -36354 42728
rect -36318 42692 -36276 42728
rect -36478 42674 -36276 42692
<< ndiffc >>
rect -37074 44950 -37038 44986
rect -37074 44806 -37038 44842
rect -37268 44672 -37234 44708
rect -37194 44672 -37160 44708
rect -37126 44672 -37092 44708
rect -37056 44672 -37020 44708
rect -37268 44528 -37234 44564
rect -37194 44528 -37160 44564
rect -37126 44528 -37092 44564
rect -37058 44528 -37022 44564
rect -37552 44256 -37518 44292
rect -37478 44256 -37444 44292
rect -37398 44256 -37364 44292
rect -37074 44256 -37038 44292
rect -37552 44112 -37516 44148
rect -37476 44112 -37440 44148
rect -37398 44114 -37364 44150
rect -37074 44112 -37038 44148
rect -37552 43984 -37518 44020
rect -37478 43984 -37444 44020
rect -37398 43984 -37364 44020
rect -37074 43984 -37038 44020
rect -37552 43840 -37516 43876
rect -37476 43840 -37440 43876
rect -37398 43842 -37364 43878
rect -37074 43840 -37038 43876
rect -37552 43712 -37518 43748
rect -37478 43712 -37444 43748
rect -37398 43712 -37364 43748
rect -37074 43712 -37038 43748
rect -37552 43568 -37516 43604
rect -37476 43568 -37440 43604
rect -37398 43570 -37364 43606
rect -37074 43568 -37038 43604
rect -37552 43440 -37518 43476
rect -37478 43440 -37444 43476
rect -37398 43440 -37364 43476
rect -37076 43440 -37040 43476
rect -37552 43296 -37516 43332
rect -37476 43296 -37440 43332
rect -37398 43298 -37364 43334
rect -37076 43296 -37040 43332
rect -37552 43168 -37518 43204
rect -37478 43168 -37444 43204
rect -37398 43168 -37364 43204
rect -37076 43168 -37040 43204
rect -37552 43024 -37516 43060
rect -37476 43024 -37440 43060
rect -37398 43026 -37364 43062
rect -37076 43024 -37040 43060
rect -37482 42838 -37448 42874
rect -37398 42838 -37364 42874
rect -37480 42694 -37444 42730
rect -37398 42694 -37362 42730
<< pdiffc >>
rect -36758 44950 -36722 44986
rect -36686 44950 -36650 44986
rect -36616 44950 -36580 44986
rect -36758 44806 -36722 44842
rect -36688 44806 -36652 44842
rect -36618 44806 -36582 44842
rect -36758 44672 -36722 44708
rect -36688 44674 -36652 44710
rect -36618 44674 -36582 44710
rect -36548 44674 -36512 44710
rect -36478 44674 -36442 44710
rect -36408 44674 -36372 44710
rect -36338 44674 -36302 44710
rect -36268 44674 -36232 44710
rect -36758 44528 -36722 44564
rect -36688 44528 -36652 44564
rect -36618 44528 -36582 44564
rect -36548 44528 -36512 44564
rect -36478 44528 -36442 44564
rect -36408 44528 -36372 44564
rect -36338 44528 -36302 44564
rect -36268 44528 -36232 44564
rect -36758 44256 -36722 44292
rect -36436 44258 -36402 44294
rect -36356 44258 -36322 44294
rect -36282 44258 -36248 44294
rect -36758 44112 -36722 44148
rect -36436 44116 -36402 44152
rect -36360 44114 -36324 44150
rect -36284 44114 -36248 44150
rect -36758 43984 -36722 44020
rect -36436 43986 -36402 44022
rect -36356 43986 -36322 44022
rect -36282 43986 -36248 44022
rect -36758 43840 -36722 43876
rect -36436 43844 -36402 43880
rect -36360 43842 -36324 43878
rect -36284 43842 -36248 43878
rect -36758 43712 -36722 43748
rect -36436 43714 -36402 43750
rect -36356 43714 -36322 43750
rect -36282 43714 -36248 43750
rect -36758 43568 -36722 43604
rect -36436 43572 -36402 43608
rect -36360 43570 -36324 43606
rect -36284 43570 -36248 43606
rect -36760 43440 -36724 43476
rect -36436 43442 -36402 43478
rect -36356 43442 -36322 43478
rect -36282 43442 -36248 43478
rect -36760 43296 -36724 43332
rect -36436 43300 -36402 43336
rect -36360 43298 -36324 43334
rect -36284 43298 -36248 43334
rect -36760 43168 -36724 43204
rect -36436 43170 -36402 43206
rect -36356 43170 -36322 43206
rect -36282 43170 -36248 43206
rect -36760 43024 -36724 43060
rect -36436 43028 -36402 43064
rect -36360 43026 -36324 43062
rect -36284 43026 -36248 43062
rect -36446 42836 -36410 42872
rect -36376 42838 -36340 42874
rect -36436 42692 -36400 42728
rect -36354 42692 -36318 42728
<< psubdiff >>
rect -37722 44722 -37686 44746
rect -37722 44662 -37686 44686
rect -37722 44446 -37686 44470
rect -37722 44386 -37686 44410
rect -37722 44104 -37686 44128
rect -37722 44044 -37686 44068
rect -37722 43830 -37686 43854
rect -37722 43770 -37686 43794
rect -37722 43558 -37686 43582
rect -37722 43498 -37686 43522
rect -37722 43288 -37686 43312
rect -37722 43228 -37686 43252
rect -37722 42966 -37686 42990
rect -37722 42906 -37686 42930
<< nsubdiff >>
rect -36116 44708 -36080 44732
rect -36116 44648 -36080 44672
rect -36116 44450 -36080 44474
rect -36116 44390 -36080 44414
rect -36116 44142 -36080 44166
rect -36116 44082 -36080 44106
rect -36116 43872 -36080 43896
rect -36116 43812 -36080 43836
rect -36116 43614 -36080 43638
rect -36116 43554 -36080 43578
rect -36124 43338 -36074 43372
rect -36124 43302 -36114 43338
rect -36078 43302 -36074 43338
rect -36124 43274 -36074 43302
rect -36114 42986 -36078 43010
rect -36114 42926 -36078 42950
<< psubdiffcont >>
rect -37722 44686 -37686 44722
rect -37722 44410 -37686 44446
rect -37722 44068 -37686 44104
rect -37722 43794 -37686 43830
rect -37722 43522 -37686 43558
rect -37722 43252 -37686 43288
rect -37722 42930 -37686 42966
<< nsubdiffcont >>
rect -36116 44672 -36080 44708
rect -36116 44414 -36080 44450
rect -36116 44106 -36080 44142
rect -36116 43836 -36080 43872
rect -36116 43578 -36080 43614
rect -36114 43302 -36078 43338
rect -36114 42950 -36078 42986
<< poly >>
rect -37160 44878 -37134 44914
rect -37004 44890 -36790 44914
rect -37004 44878 -36910 44890
rect -36926 44854 -36910 44878
rect -36874 44878 -36790 44890
rect -36532 44878 -36506 44914
rect -36874 44854 -36858 44878
rect -36926 44840 -36858 44854
rect -36914 44830 -36870 44840
rect -37318 44600 -37292 44636
rect -37004 44612 -36790 44636
rect -37004 44600 -36910 44612
rect -36926 44576 -36910 44600
rect -36874 44600 -36790 44612
rect -36214 44600 -36188 44636
rect -36874 44576 -36858 44600
rect -36926 44562 -36858 44576
rect -36914 44552 -36870 44562
rect -37278 44256 -37234 44266
rect -37290 44242 -37222 44256
rect -37290 44220 -37274 44242
rect -37608 44184 -37582 44220
rect -37324 44206 -37274 44220
rect -37238 44206 -37222 44242
rect -36566 44258 -36522 44268
rect -36578 44244 -36510 44258
rect -37324 44184 -37222 44206
rect -37142 44184 -37106 44220
rect -37006 44196 -36790 44220
rect -37006 44184 -36910 44196
rect -36926 44160 -36910 44184
rect -36874 44184 -36790 44196
rect -36690 44184 -36654 44220
rect -36578 44208 -36562 44244
rect -36526 44222 -36510 44244
rect -36526 44208 -36478 44222
rect -36578 44186 -36478 44208
rect -36218 44186 -36192 44222
rect -36874 44160 -36858 44184
rect -36926 44146 -36858 44160
rect -36914 44136 -36870 44146
rect -37278 43984 -37234 43994
rect -37290 43970 -37222 43984
rect -37290 43948 -37274 43970
rect -37608 43912 -37582 43948
rect -37324 43934 -37274 43948
rect -37238 43934 -37222 43970
rect -36566 43986 -36522 43996
rect -36578 43972 -36510 43986
rect -37324 43912 -37222 43934
rect -37142 43912 -37106 43948
rect -37006 43924 -36790 43948
rect -37006 43912 -36910 43924
rect -36926 43888 -36910 43912
rect -36874 43912 -36790 43924
rect -36690 43912 -36654 43948
rect -36578 43936 -36562 43972
rect -36526 43950 -36510 43972
rect -36526 43936 -36478 43950
rect -36578 43914 -36478 43936
rect -36218 43914 -36192 43950
rect -36874 43888 -36858 43912
rect -36926 43874 -36858 43888
rect -36914 43864 -36870 43874
rect -37278 43712 -37234 43722
rect -37290 43698 -37222 43712
rect -37290 43676 -37274 43698
rect -37608 43640 -37582 43676
rect -37324 43662 -37274 43676
rect -37238 43662 -37222 43698
rect -36566 43714 -36522 43724
rect -36578 43700 -36510 43714
rect -37324 43640 -37222 43662
rect -37142 43640 -37106 43676
rect -37006 43652 -36790 43676
rect -37006 43640 -36910 43652
rect -36926 43616 -36910 43640
rect -36874 43640 -36790 43652
rect -36690 43640 -36654 43676
rect -36578 43664 -36562 43700
rect -36526 43678 -36510 43700
rect -36526 43664 -36478 43678
rect -36578 43642 -36478 43664
rect -36218 43642 -36192 43678
rect -36874 43616 -36858 43640
rect -36926 43602 -36858 43616
rect -36914 43592 -36870 43602
rect -37278 43440 -37234 43450
rect -37290 43426 -37222 43440
rect -37290 43404 -37274 43426
rect -37608 43368 -37582 43404
rect -37324 43390 -37274 43404
rect -37238 43390 -37222 43426
rect -36566 43442 -36522 43452
rect -36578 43428 -36510 43442
rect -37324 43368 -37222 43390
rect -37144 43368 -37108 43404
rect -37008 43380 -36792 43404
rect -37008 43368 -36912 43380
rect -36928 43344 -36912 43368
rect -36876 43368 -36792 43380
rect -36692 43368 -36656 43404
rect -36578 43392 -36562 43428
rect -36526 43406 -36510 43428
rect -36526 43392 -36478 43406
rect -36578 43370 -36478 43392
rect -36218 43370 -36192 43406
rect -36876 43344 -36860 43368
rect -36928 43330 -36860 43344
rect -36916 43320 -36872 43330
rect -37278 43168 -37234 43178
rect -37290 43154 -37222 43168
rect -37290 43132 -37274 43154
rect -37608 43096 -37582 43132
rect -37324 43118 -37274 43132
rect -37238 43118 -37222 43154
rect -36566 43170 -36522 43180
rect -36578 43156 -36510 43170
rect -37324 43096 -37222 43118
rect -37144 43096 -37108 43132
rect -37008 43108 -36792 43132
rect -37008 43096 -36912 43108
rect -36928 43072 -36912 43096
rect -36876 43096 -36792 43108
rect -36692 43096 -36656 43132
rect -36578 43120 -36562 43156
rect -36526 43134 -36510 43156
rect -36526 43120 -36478 43134
rect -36578 43098 -36478 43120
rect -36218 43098 -36192 43134
rect -36876 43072 -36860 43096
rect -36928 43058 -36860 43072
rect -36916 43048 -36872 43058
rect -37278 42838 -37234 42848
rect -37290 42824 -37222 42838
rect -36566 42836 -36522 42846
rect -37290 42802 -37274 42824
rect -37550 42766 -37524 42802
rect -37322 42788 -37274 42802
rect -37238 42788 -37222 42824
rect -37322 42766 -37222 42788
rect -36578 42822 -36510 42836
rect -36578 42786 -36562 42822
rect -36526 42800 -36510 42822
rect -36526 42786 -36478 42800
rect -36578 42764 -36478 42786
rect -36276 42764 -36250 42800
<< polycont >>
rect -36910 44854 -36874 44890
rect -36910 44576 -36874 44612
rect -37274 44206 -37238 44242
rect -36910 44160 -36874 44196
rect -36562 44208 -36526 44244
rect -37274 43934 -37238 43970
rect -36910 43888 -36874 43924
rect -36562 43936 -36526 43972
rect -37274 43662 -37238 43698
rect -36910 43616 -36874 43652
rect -36562 43664 -36526 43700
rect -37274 43390 -37238 43426
rect -36912 43344 -36876 43380
rect -36562 43392 -36526 43428
rect -37274 43118 -37238 43154
rect -36912 43072 -36876 43108
rect -36562 43120 -36526 43156
rect -37274 42788 -37238 42824
rect -36562 42786 -36526 42822
<< locali >>
rect -37090 44990 -37006 45002
rect -36910 44990 -36874 45030
rect -36790 44990 -36540 45002
rect -37090 44986 -36540 44990
rect -37090 44950 -37074 44986
rect -37038 44950 -36758 44986
rect -36722 44950 -36686 44986
rect -36650 44950 -36616 44986
rect -36580 44950 -36540 44986
rect -37090 44946 -36540 44950
rect -37090 44934 -37006 44946
rect -36790 44934 -36540 44946
rect -37744 44856 -37666 44900
rect -36926 44890 -36858 44900
rect -37094 44856 -37022 44858
rect -37744 44844 -37022 44856
rect -36926 44854 -36910 44890
rect -36874 44854 -36858 44890
rect -36138 44858 -36064 44872
rect -36926 44846 -36858 44854
rect -37744 44808 -37722 44844
rect -37686 44842 -37022 44844
rect -37686 44808 -37074 44842
rect -37744 44806 -37074 44808
rect -37038 44806 -37022 44842
rect -37744 44794 -37022 44806
rect -37744 44722 -37666 44794
rect -37094 44790 -37022 44794
rect -37744 44686 -37722 44722
rect -37686 44686 -37666 44722
rect -37744 44580 -37666 44686
rect -37276 44712 -37006 44724
rect -36910 44712 -36874 44846
rect -36778 44842 -36064 44858
rect -36778 44806 -36758 44842
rect -36722 44806 -36688 44842
rect -36652 44806 -36618 44842
rect -36582 44806 -36118 44842
rect -36082 44806 -36064 44842
rect -36778 44790 -36064 44806
rect -36790 44720 -36708 44724
rect -36790 44712 -36216 44720
rect -37276 44710 -36216 44712
rect -37276 44708 -36688 44710
rect -37276 44672 -37268 44708
rect -37234 44672 -37194 44708
rect -37160 44672 -37126 44708
rect -37092 44672 -37056 44708
rect -37020 44672 -36758 44708
rect -36722 44674 -36688 44708
rect -36652 44674 -36618 44710
rect -36582 44674 -36548 44710
rect -36512 44674 -36478 44710
rect -36442 44674 -36408 44710
rect -36372 44674 -36338 44710
rect -36302 44674 -36268 44710
rect -36232 44674 -36216 44710
rect -36722 44672 -36216 44674
rect -37276 44668 -36216 44672
rect -37276 44658 -37006 44668
rect -37268 44656 -37006 44658
rect -36790 44656 -36216 44668
rect -36138 44708 -36064 44790
rect -36138 44672 -36116 44708
rect -36080 44672 -36064 44708
rect -36926 44612 -36858 44622
rect -37744 44564 -37008 44580
rect -36926 44576 -36910 44612
rect -36874 44576 -36858 44612
rect -36138 44582 -36064 44672
rect -36236 44580 -36064 44582
rect -36926 44568 -36858 44576
rect -37744 44558 -37268 44564
rect -37744 44522 -37722 44558
rect -37686 44528 -37268 44558
rect -37234 44528 -37194 44564
rect -37160 44528 -37126 44564
rect -37092 44528 -37058 44564
rect -37022 44528 -37008 44564
rect -37686 44522 -37008 44528
rect -37744 44514 -37008 44522
rect -37744 44512 -37022 44514
rect -37744 44446 -37666 44512
rect -37744 44410 -37722 44446
rect -37686 44410 -37666 44446
rect -37744 44306 -37666 44410
rect -36910 44364 -36874 44568
rect -36778 44566 -36064 44580
rect -36778 44564 -36118 44566
rect -36778 44528 -36758 44564
rect -36722 44528 -36688 44564
rect -36652 44528 -36618 44564
rect -36582 44528 -36548 44564
rect -36512 44528 -36478 44564
rect -36442 44528 -36408 44564
rect -36372 44528 -36338 44564
rect -36302 44528 -36268 44564
rect -36232 44530 -36118 44564
rect -36082 44530 -36064 44566
rect -36232 44528 -36064 44530
rect -36778 44514 -36064 44528
rect -36778 44512 -36222 44514
rect -36138 44450 -36064 44514
rect -36138 44414 -36116 44450
rect -36080 44414 -36064 44450
rect -37582 44306 -37338 44308
rect -37744 44292 -37338 44306
rect -37744 44290 -37552 44292
rect -37744 44254 -37722 44290
rect -37686 44256 -37552 44290
rect -37518 44256 -37478 44292
rect -37444 44256 -37398 44292
rect -37364 44256 -37338 44292
rect -37686 44254 -37338 44256
rect -37744 44242 -37338 44254
rect -37274 44250 -37238 44284
rect -37090 44296 -37006 44308
rect -36910 44296 -36874 44322
rect -36790 44296 -36708 44308
rect -37090 44292 -36708 44296
rect -37090 44256 -37074 44292
rect -37038 44256 -36758 44292
rect -36722 44256 -36708 44292
rect -37090 44252 -36708 44256
rect -36138 44312 -36064 44414
rect -36222 44310 -36064 44312
rect -36562 44252 -36526 44286
rect -36462 44306 -36064 44310
rect -36462 44296 -36062 44306
rect -36462 44294 -36118 44296
rect -36462 44258 -36436 44294
rect -36402 44258 -36356 44294
rect -36322 44258 -36282 44294
rect -36248 44260 -36118 44294
rect -36082 44260 -36062 44296
rect -36248 44258 -36062 44260
rect -37744 44104 -37666 44242
rect -37582 44240 -37338 44242
rect -37290 44242 -37222 44250
rect -37290 44206 -37274 44242
rect -37238 44206 -37222 44242
rect -37090 44240 -37006 44252
rect -36790 44240 -36708 44252
rect -36578 44244 -36510 44252
rect -36578 44208 -36562 44244
rect -36526 44208 -36510 44244
rect -36462 44244 -36062 44258
rect -36462 44242 -36218 44244
rect -37290 44196 -37222 44206
rect -36926 44196 -36858 44206
rect -36578 44198 -36510 44208
rect -37744 44068 -37722 44104
rect -37686 44068 -37666 44104
rect -37582 44154 -37324 44166
rect -37582 44152 -37322 44154
rect -37094 44152 -37022 44164
rect -36926 44160 -36910 44196
rect -36874 44160 -36858 44196
rect -36926 44152 -36858 44160
rect -36778 44154 -36706 44164
rect -36476 44156 -36218 44168
rect -36478 44154 -36218 44156
rect -36778 44152 -36218 44154
rect -37582 44150 -37022 44152
rect -37582 44148 -37398 44150
rect -37582 44112 -37552 44148
rect -37516 44112 -37476 44148
rect -37440 44114 -37398 44148
rect -37364 44148 -37022 44150
rect -37364 44114 -37074 44148
rect -37440 44112 -37074 44114
rect -37038 44112 -37022 44148
rect -37582 44106 -37022 44112
rect -37582 44096 -37324 44106
rect -37094 44096 -37022 44106
rect -37744 44034 -37666 44068
rect -37582 44034 -37338 44036
rect -37744 44020 -37338 44034
rect -37744 43984 -37552 44020
rect -37518 43984 -37478 44020
rect -37444 43984 -37398 44020
rect -37364 43984 -37338 44020
rect -37744 43970 -37338 43984
rect -37274 43978 -37238 44012
rect -37090 44024 -37006 44036
rect -36910 44024 -36874 44152
rect -36778 44148 -36436 44152
rect -36778 44112 -36758 44148
rect -36722 44116 -36436 44148
rect -36402 44150 -36218 44152
rect -36402 44116 -36360 44150
rect -36722 44114 -36360 44116
rect -36324 44114 -36284 44150
rect -36248 44114 -36218 44150
rect -36722 44112 -36218 44114
rect -36778 44108 -36218 44112
rect -36778 44096 -36706 44108
rect -36476 44098 -36218 44108
rect -36138 44142 -36062 44244
rect -36138 44106 -36116 44142
rect -36080 44106 -36062 44142
rect -36790 44024 -36708 44036
rect -37090 44020 -36708 44024
rect -37090 43984 -37074 44020
rect -37038 43984 -36758 44020
rect -36722 43984 -36708 44020
rect -37090 43980 -36708 43984
rect -36138 44040 -36062 44106
rect -36220 44038 -36062 44040
rect -36562 43980 -36526 44014
rect -36462 44022 -36062 44038
rect -36462 43986 -36436 44022
rect -36402 43986 -36356 44022
rect -36322 43986 -36282 44022
rect -36248 43986 -36116 44022
rect -36080 43986 -36062 44022
rect -37744 43934 -37722 43970
rect -37686 43934 -37666 43970
rect -37582 43968 -37338 43970
rect -37290 43970 -37222 43978
rect -37744 43830 -37666 43934
rect -37290 43934 -37274 43970
rect -37238 43934 -37222 43970
rect -37090 43968 -37006 43980
rect -36790 43968 -36708 43980
rect -36578 43972 -36510 43980
rect -36578 43936 -36562 43972
rect -36526 43936 -36510 43972
rect -36462 43972 -36062 43986
rect -36462 43970 -36218 43972
rect -37290 43924 -37222 43934
rect -36926 43924 -36858 43934
rect -36578 43926 -36510 43936
rect -37744 43794 -37722 43830
rect -37686 43794 -37666 43830
rect -37582 43882 -37324 43894
rect -37582 43880 -37322 43882
rect -37094 43880 -37022 43892
rect -36926 43888 -36910 43924
rect -36874 43888 -36858 43924
rect -36926 43880 -36858 43888
rect -36778 43882 -36706 43892
rect -36476 43884 -36218 43896
rect -36478 43882 -36218 43884
rect -36778 43880 -36218 43882
rect -37582 43878 -37022 43880
rect -37582 43876 -37398 43878
rect -37582 43840 -37552 43876
rect -37516 43840 -37476 43876
rect -37440 43842 -37398 43876
rect -37364 43876 -37022 43878
rect -37364 43842 -37074 43876
rect -37440 43840 -37074 43842
rect -37038 43840 -37022 43876
rect -37582 43834 -37022 43840
rect -37582 43824 -37324 43834
rect -37094 43824 -37022 43834
rect -37744 43764 -37666 43794
rect -37744 43748 -37338 43764
rect -37744 43712 -37552 43748
rect -37518 43712 -37478 43748
rect -37444 43712 -37398 43748
rect -37364 43712 -37338 43748
rect -37744 43700 -37338 43712
rect -37274 43706 -37238 43740
rect -37090 43752 -37006 43764
rect -36910 43752 -36874 43880
rect -36778 43876 -36436 43880
rect -36778 43840 -36758 43876
rect -36722 43844 -36436 43876
rect -36402 43878 -36218 43880
rect -36402 43844 -36360 43878
rect -36722 43842 -36360 43844
rect -36324 43842 -36284 43878
rect -36248 43842 -36218 43878
rect -36722 43840 -36218 43842
rect -36778 43836 -36218 43840
rect -36778 43824 -36706 43836
rect -36476 43826 -36218 43836
rect -36138 43872 -36062 43972
rect -36138 43836 -36116 43872
rect -36080 43836 -36062 43872
rect -36790 43752 -36708 43764
rect -37090 43748 -36708 43752
rect -37090 43712 -37074 43748
rect -37038 43712 -36758 43748
rect -36722 43712 -36708 43748
rect -37090 43708 -36708 43712
rect -36138 43766 -36062 43836
rect -36562 43708 -36526 43742
rect -36462 43750 -36062 43766
rect -36462 43714 -36436 43750
rect -36402 43714 -36356 43750
rect -36322 43714 -36282 43750
rect -36248 43714 -36114 43750
rect -36078 43714 -36062 43750
rect -37744 43694 -37666 43700
rect -37582 43696 -37338 43700
rect -37290 43698 -37222 43706
rect -37744 43658 -37722 43694
rect -37686 43658 -37666 43694
rect -37744 43558 -37666 43658
rect -37290 43662 -37274 43698
rect -37238 43662 -37222 43698
rect -37090 43696 -37006 43708
rect -36790 43696 -36708 43708
rect -36578 43700 -36510 43708
rect -36578 43664 -36562 43700
rect -36526 43664 -36510 43700
rect -36462 43698 -36062 43714
rect -37290 43652 -37222 43662
rect -36926 43652 -36858 43662
rect -36578 43654 -36510 43664
rect -37744 43522 -37722 43558
rect -37686 43522 -37666 43558
rect -37582 43610 -37324 43622
rect -37582 43608 -37322 43610
rect -37094 43608 -37022 43620
rect -36926 43616 -36910 43652
rect -36874 43616 -36858 43652
rect -36926 43608 -36858 43616
rect -36778 43610 -36706 43620
rect -36476 43612 -36218 43624
rect -36478 43610 -36218 43612
rect -36778 43608 -36218 43610
rect -37582 43606 -37022 43608
rect -37582 43604 -37398 43606
rect -37582 43568 -37552 43604
rect -37516 43568 -37476 43604
rect -37440 43570 -37398 43604
rect -37364 43604 -37022 43606
rect -37364 43570 -37074 43604
rect -37440 43568 -37074 43570
rect -37038 43568 -37022 43604
rect -37582 43562 -37022 43568
rect -37582 43552 -37324 43562
rect -37094 43552 -37022 43562
rect -36910 43560 -36874 43608
rect -37744 43490 -37666 43522
rect -36912 43532 -36874 43560
rect -36778 43604 -36436 43608
rect -36778 43568 -36758 43604
rect -36722 43572 -36436 43604
rect -36402 43606 -36218 43608
rect -36402 43572 -36360 43606
rect -36722 43570 -36360 43572
rect -36324 43570 -36284 43606
rect -36248 43570 -36218 43606
rect -36722 43568 -36218 43570
rect -36778 43564 -36218 43568
rect -36778 43552 -36706 43564
rect -36476 43554 -36218 43564
rect -36138 43614 -36062 43698
rect -36138 43578 -36116 43614
rect -36080 43578 -36062 43614
rect -37582 43490 -37338 43492
rect -37744 43476 -37338 43490
rect -37744 43440 -37552 43476
rect -37518 43440 -37478 43476
rect -37444 43440 -37398 43476
rect -37364 43440 -37338 43476
rect -37744 43426 -37338 43440
rect -37274 43434 -37238 43468
rect -37092 43480 -37008 43492
rect -36912 43480 -36876 43532
rect -36792 43480 -36710 43492
rect -37092 43476 -36710 43480
rect -37092 43440 -37076 43476
rect -37040 43440 -36760 43476
rect -36724 43440 -36710 43476
rect -37092 43436 -36710 43440
rect -36138 43494 -36062 43578
rect -36562 43436 -36526 43470
rect -36462 43480 -36062 43494
rect -36462 43478 -36114 43480
rect -36462 43442 -36436 43478
rect -36402 43442 -36356 43478
rect -36322 43442 -36282 43478
rect -36248 43444 -36114 43478
rect -36078 43444 -36062 43480
rect -36248 43442 -36062 43444
rect -37744 43422 -37666 43426
rect -37582 43424 -37338 43426
rect -37290 43426 -37222 43434
rect -37744 43386 -37722 43422
rect -37686 43386 -37666 43422
rect -37744 43288 -37666 43386
rect -37290 43390 -37274 43426
rect -37238 43390 -37222 43426
rect -37092 43424 -37008 43436
rect -36792 43424 -36710 43436
rect -36578 43428 -36510 43436
rect -36578 43392 -36562 43428
rect -36526 43392 -36510 43428
rect -36462 43426 -36062 43442
rect -37290 43380 -37222 43390
rect -36928 43380 -36860 43390
rect -36578 43382 -36510 43392
rect -37744 43252 -37722 43288
rect -37686 43252 -37666 43288
rect -37582 43338 -37324 43350
rect -37582 43336 -37322 43338
rect -37096 43336 -37024 43348
rect -36928 43344 -36912 43380
rect -36876 43344 -36860 43380
rect -36928 43336 -36860 43344
rect -36780 43338 -36708 43348
rect -36476 43340 -36218 43352
rect -36478 43338 -36218 43340
rect -36780 43336 -36218 43338
rect -37582 43334 -37024 43336
rect -37582 43332 -37398 43334
rect -37582 43296 -37552 43332
rect -37516 43296 -37476 43332
rect -37440 43298 -37398 43332
rect -37364 43332 -37024 43334
rect -37364 43298 -37076 43332
rect -37440 43296 -37076 43298
rect -37040 43296 -37024 43332
rect -37582 43290 -37024 43296
rect -37582 43280 -37324 43290
rect -37096 43280 -37024 43290
rect -37744 43218 -37666 43252
rect -37582 43218 -37338 43220
rect -37744 43204 -37338 43218
rect -37744 43168 -37552 43204
rect -37518 43168 -37478 43204
rect -37444 43168 -37398 43204
rect -37364 43168 -37338 43204
rect -37744 43154 -37338 43168
rect -37274 43162 -37238 43196
rect -37092 43208 -37008 43220
rect -36912 43208 -36876 43336
rect -36780 43332 -36436 43336
rect -36780 43296 -36760 43332
rect -36724 43300 -36436 43332
rect -36402 43334 -36218 43336
rect -36402 43300 -36360 43334
rect -36724 43298 -36360 43300
rect -36324 43298 -36284 43334
rect -36248 43298 -36218 43334
rect -36724 43296 -36218 43298
rect -36780 43292 -36218 43296
rect -36780 43280 -36708 43292
rect -36476 43282 -36218 43292
rect -36138 43338 -36062 43426
rect -36138 43302 -36114 43338
rect -36078 43302 -36062 43338
rect -36792 43208 -36710 43220
rect -37092 43204 -36710 43208
rect -37092 43168 -37076 43204
rect -37040 43168 -36760 43204
rect -36724 43168 -36710 43204
rect -37092 43164 -36710 43168
rect -36138 43224 -36062 43302
rect -36218 43222 -36062 43224
rect -36562 43164 -36526 43198
rect -36462 43208 -36062 43222
rect -36462 43206 -36114 43208
rect -36462 43170 -36436 43206
rect -36402 43170 -36356 43206
rect -36322 43170 -36282 43206
rect -36248 43172 -36114 43206
rect -36078 43172 -36062 43208
rect -36248 43170 -36062 43172
rect -37744 43110 -37666 43154
rect -37582 43152 -37338 43154
rect -37290 43154 -37222 43162
rect -37744 43074 -37722 43110
rect -37686 43074 -37666 43110
rect -37290 43118 -37274 43154
rect -37238 43118 -37222 43154
rect -37092 43152 -37008 43164
rect -36792 43152 -36710 43164
rect -36578 43156 -36510 43164
rect -36578 43120 -36562 43156
rect -36526 43120 -36510 43156
rect -36462 43156 -36062 43170
rect -36462 43154 -36218 43156
rect -36138 43154 -36062 43156
rect -37290 43108 -37222 43118
rect -36928 43108 -36860 43118
rect -36578 43110 -36510 43120
rect -37744 42966 -37666 43074
rect -37582 43066 -37324 43078
rect -37582 43064 -37322 43066
rect -37096 43064 -37024 43076
rect -36928 43072 -36912 43108
rect -36876 43072 -36860 43108
rect -36928 43064 -36860 43072
rect -36780 43066 -36708 43076
rect -36476 43068 -36218 43080
rect -36478 43066 -36218 43068
rect -36780 43064 -36218 43066
rect -37582 43062 -37024 43064
rect -37582 43060 -37398 43062
rect -37582 43024 -37552 43060
rect -37516 43024 -37476 43060
rect -37440 43026 -37398 43060
rect -37364 43060 -37024 43062
rect -37364 43026 -37076 43060
rect -37440 43024 -37076 43026
rect -37040 43024 -37024 43060
rect -37582 43018 -37024 43024
rect -37582 43008 -37324 43018
rect -37096 43008 -37024 43018
rect -36912 43030 -36876 43064
rect -36780 43060 -36436 43064
rect -36780 43024 -36760 43060
rect -36724 43028 -36436 43060
rect -36402 43062 -36218 43064
rect -36402 43028 -36360 43062
rect -36724 43026 -36360 43028
rect -36324 43026 -36284 43062
rect -36248 43026 -36218 43062
rect -36724 43024 -36218 43026
rect -36780 43020 -36218 43024
rect -36780 43008 -36708 43020
rect -36476 43010 -36218 43020
rect -37744 42930 -37722 42966
rect -37686 42930 -37666 42966
rect -37744 42884 -37666 42930
rect -36136 42986 -36062 43154
rect -36136 42950 -36114 42986
rect -36078 42950 -36062 42986
rect -37524 42884 -37342 42890
rect -37744 42874 -37342 42884
rect -37744 42872 -37482 42874
rect -37744 42836 -37722 42872
rect -37686 42838 -37482 42872
rect -37448 42838 -37398 42874
rect -37364 42838 -37342 42874
rect -37686 42836 -37342 42838
rect -37744 42830 -37342 42836
rect -37274 42832 -37238 42866
rect -36136 42884 -36062 42950
rect -37744 42770 -37666 42830
rect -37524 42822 -37342 42830
rect -37290 42824 -37222 42832
rect -36562 42830 -36526 42864
rect -36466 42874 -36062 42884
rect -36466 42872 -36376 42874
rect -36466 42836 -36446 42872
rect -36410 42838 -36376 42872
rect -36340 42868 -36062 42874
rect -36340 42838 -36114 42868
rect -36410 42836 -36114 42838
rect -36466 42832 -36114 42836
rect -36078 42832 -36062 42868
rect -37290 42788 -37274 42824
rect -37238 42788 -37222 42824
rect -37290 42778 -37222 42788
rect -36578 42822 -36510 42830
rect -36578 42786 -36562 42822
rect -36526 42786 -36510 42822
rect -36466 42820 -36062 42832
rect -36578 42776 -36510 42786
rect -37524 42736 -37342 42748
rect -36572 42740 -36522 42776
rect -36474 42740 -36294 42744
rect -36572 42736 -36294 42740
rect -37524 42730 -36294 42736
rect -37524 42694 -37480 42730
rect -37444 42694 -37398 42730
rect -37362 42728 -36294 42730
rect -37362 42694 -36436 42728
rect -37524 42692 -36436 42694
rect -36400 42692 -36354 42728
rect -36318 42692 -36294 42728
rect -37524 42684 -36294 42692
rect -37524 42678 -37342 42684
rect -36572 42682 -36294 42684
rect -36478 42676 -36294 42682
rect -36136 42586 -36062 42820
rect -36136 42396 -36064 42586
rect -36134 42230 -36064 42396
rect -36134 42192 -36118 42230
rect -36080 42192 -36064 42230
rect -36134 42182 -36064 42192
<< viali >>
rect -36910 45030 -36874 45066
rect -37722 44808 -37686 44844
rect -36118 44806 -36082 44842
rect -37722 44522 -37686 44558
rect -36118 44530 -36082 44566
rect -36910 44322 -36874 44364
rect -37722 44254 -37686 44290
rect -37274 44284 -37238 44322
rect -36562 44286 -36526 44324
rect -36118 44260 -36082 44296
rect -37274 44012 -37238 44050
rect -36562 44014 -36526 44052
rect -36116 43986 -36080 44022
rect -37722 43934 -37686 43970
rect -37274 43740 -37238 43778
rect -36562 43742 -36526 43780
rect -36114 43714 -36078 43750
rect -37722 43658 -37686 43694
rect -37274 43468 -37238 43506
rect -36562 43470 -36526 43508
rect -36114 43444 -36078 43480
rect -37722 43386 -37686 43422
rect -37274 43196 -37238 43234
rect -36562 43198 -36526 43236
rect -36114 43172 -36078 43208
rect -37722 43074 -37686 43110
rect -36912 42988 -36876 43030
rect -37722 42836 -37686 42872
rect -37274 42866 -37238 42904
rect -36562 42864 -36526 42902
rect -36114 42832 -36078 42868
rect -36118 42192 -36080 42230
<< metal1 >>
rect -36926 45220 -36856 45300
rect -36930 45210 -36852 45220
rect -36930 45154 -36918 45210
rect -36862 45154 -36852 45210
rect -36930 45134 -36852 45154
rect -36922 45066 -36864 45134
rect -37740 44982 -37670 45062
rect -36922 45030 -36910 45066
rect -36874 45030 -36864 45066
rect -36922 45000 -36864 45030
rect -37744 44972 -37666 44982
rect -37744 44916 -37732 44972
rect -37676 44916 -37666 44972
rect -37744 44900 -37666 44916
rect -37746 44896 -37666 44900
rect -37746 44844 -37664 44896
rect -37746 44808 -37722 44844
rect -37686 44808 -37664 44844
rect -37746 44558 -37664 44808
rect -37746 44522 -37722 44558
rect -37686 44522 -37664 44558
rect -37746 44290 -37664 44522
rect -36134 44842 -36062 44870
rect -36134 44806 -36118 44842
rect -36082 44806 -36062 44842
rect -36134 44566 -36062 44806
rect -36134 44530 -36118 44566
rect -36082 44530 -36062 44566
rect -36922 44364 -36864 44376
rect -37746 44254 -37722 44290
rect -37686 44254 -37664 44290
rect -37746 43970 -37664 44254
rect -37746 43934 -37722 43970
rect -37686 43934 -37664 43970
rect -37746 43694 -37664 43934
rect -37746 43658 -37722 43694
rect -37686 43658 -37664 43694
rect -37746 43422 -37664 43658
rect -37746 43386 -37722 43422
rect -37686 43386 -37664 43422
rect -37746 43110 -37664 43386
rect -37746 43074 -37722 43110
rect -37686 43074 -37664 43110
rect -37746 42872 -37664 43074
rect -37746 42836 -37722 42872
rect -37686 42836 -37664 42872
rect -37746 42768 -37664 42836
rect -37284 44322 -37226 44336
rect -37284 44284 -37274 44322
rect -37238 44284 -37226 44322
rect -37284 44050 -37226 44284
rect -37284 44012 -37274 44050
rect -37238 44012 -37226 44050
rect -37284 43778 -37226 44012
rect -37284 43740 -37274 43778
rect -37238 43740 -37226 43778
rect -37284 43506 -37226 43740
rect -37284 43468 -37274 43506
rect -37238 43468 -37226 43506
rect -37284 43234 -37226 43468
rect -37284 43196 -37274 43234
rect -37238 43196 -37226 43234
rect -37284 42904 -37226 43196
rect -36922 44322 -36910 44364
rect -36874 44322 -36864 44364
rect -36922 43030 -36864 44322
rect -36922 42988 -36912 43030
rect -36876 42988 -36864 43030
rect -36922 42965 -36864 42988
rect -36574 44324 -36516 44338
rect -36574 44286 -36562 44324
rect -36526 44286 -36516 44324
rect -36574 44052 -36516 44286
rect -36574 44014 -36562 44052
rect -36526 44014 -36516 44052
rect -36574 43780 -36516 44014
rect -36574 43742 -36562 43780
rect -36526 43742 -36516 43780
rect -36574 43508 -36516 43742
rect -36574 43470 -36562 43508
rect -36526 43470 -36516 43508
rect -36574 43236 -36516 43470
rect -36574 43198 -36562 43236
rect -36526 43198 -36516 43236
rect -37284 42866 -37274 42904
rect -37238 42866 -37226 42904
rect -37284 42838 -37226 42866
rect -36574 42902 -36516 43198
rect -36134 44296 -36062 44530
rect -36134 44260 -36118 44296
rect -36082 44260 -36062 44296
rect -36134 44022 -36062 44260
rect -36134 43986 -36116 44022
rect -36080 43986 -36062 44022
rect -36134 43750 -36062 43986
rect -36134 43714 -36114 43750
rect -36078 43714 -36062 43750
rect -36134 43480 -36062 43714
rect -36134 43444 -36114 43480
rect -36078 43444 -36062 43480
rect -36134 43208 -36062 43444
rect -36134 43172 -36114 43208
rect -36078 43172 -36062 43208
rect -36134 43148 -36062 43172
rect -36574 42864 -36562 42902
rect -36526 42864 -36516 42902
rect -37177 42838 -36864 42841
rect -37284 42766 -36864 42838
rect -37177 42765 -36864 42766
rect -36922 42528 -36864 42765
rect -36574 42764 -36516 42864
rect -36136 42868 -36062 43148
rect -36136 42832 -36114 42868
rect -36078 42832 -36062 42868
rect -36136 42768 -36062 42832
rect -36923 42527 -36847 42528
rect -36941 42409 -36833 42527
rect -36927 42395 -36849 42409
rect -36927 42339 -36917 42395
rect -36861 42339 -36849 42395
rect -36927 42329 -36849 42339
rect -36923 42249 -36853 42329
rect -36132 42230 -36066 42246
rect -36132 42192 -36118 42230
rect -36080 42192 -36066 42230
rect -36132 42184 -36066 42192
rect -36128 42136 -36070 42184
rect -36140 42116 -36062 42136
rect -36140 42060 -36130 42116
rect -36074 42060 -36062 42116
rect -36140 42050 -36062 42060
rect -36136 41970 -36066 42050
<< via1 >>
rect -36918 45154 -36862 45210
rect -37732 44916 -37676 44972
rect -36917 42339 -36861 42395
rect -36130 42060 -36074 42116
<< metal2 >>
rect -36588 45674 -36502 45678
rect -36588 45671 -36422 45674
rect -37741 45666 -36422 45671
rect -37741 45610 -36568 45666
rect -36512 45610 -36422 45666
rect -37741 45604 -36422 45610
rect -37741 45600 -36502 45604
rect -37741 45599 -36521 45600
rect -37741 45027 -37669 45599
rect -36926 45220 -36856 45300
rect -36930 45210 -36852 45220
rect -36930 45154 -36918 45210
rect -36862 45154 -36852 45210
rect -36930 45134 -36852 45154
rect -37740 44982 -37670 45027
rect -37744 44972 -37666 44982
rect -37744 44916 -37732 44972
rect -37676 44916 -37666 44972
rect -37744 44896 -37666 44916
rect -36927 42395 -36849 42415
rect -36927 42339 -36917 42395
rect -36861 42339 -36849 42395
rect -36927 42329 -36849 42339
rect -36923 42249 -36853 42329
rect -36140 42116 -36062 42136
rect -36140 42060 -36130 42116
rect -36074 42060 -36062 42116
rect -36140 42050 -36062 42060
rect -36136 41970 -36066 42050
<< via2 >>
rect -36568 45610 -36512 45666
rect -36918 45154 -36862 45210
rect -36917 42339 -36861 42395
rect -36130 42060 -36074 42116
<< metal3 >>
rect -177846 53178 -177142 53248
rect -76328 53202 -75634 53272
rect 7950 53210 8502 53276
rect -177498 46745 -177428 53178
rect -76002 49257 -75932 53202
rect 8236 51757 8302 53210
rect 60002 53147 60548 53218
rect 8236 51704 8493 51757
rect 8237 51691 8493 51704
rect -76002 49187 -74189 49257
rect -76002 49186 -75932 49187
rect -177498 46678 -174829 46745
rect -177485 46675 -174829 46678
rect -174899 42150 -174829 46675
rect -74259 45795 -74189 49187
rect 8427 46941 8493 51691
rect -36340 46875 8493 46941
rect -74260 45725 -36856 45795
rect -36926 45220 -36856 45725
rect -36588 45674 -36502 45678
rect -36588 45671 -36405 45674
rect -36340 45671 -36274 46875
rect -36588 45666 -36274 45671
rect -36588 45610 -36568 45666
rect -36512 45610 -36274 45666
rect -36588 45605 -36274 45610
rect -36588 45604 -36405 45605
rect -36588 45600 -36502 45604
rect -36930 45210 -36852 45220
rect -36930 45154 -36918 45210
rect -36862 45154 -36852 45210
rect -36930 45134 -36852 45154
rect -36927 42395 -36849 42415
rect -36927 42339 -36917 42395
rect -36861 42339 -36849 42395
rect -36927 42329 -36849 42339
rect -36923 42150 -36853 42329
rect -174899 42080 -36853 42150
rect -36140 42116 -36062 42136
rect -36140 42060 -36130 42116
rect -36074 42060 -36062 42116
rect -36140 42050 -36062 42060
rect -36136 41985 -36066 42050
rect -36136 41299 -36065 41985
rect 60253 41299 60324 53147
rect -36136 41228 60324 41299
<< labels >>
rlabel metal3 -36455 45639 -36455 45639 1 io_analog[3]
rlabel metal3 -36891 45245 -36891 45245 1 io_analog[4]
rlabel metal3 -36889 42293 -36889 42293 1 io_analog[5]
rlabel metal3 -36103 42011 -36103 42011 1 io_analog[2]
<< end >>
