magic
tech sky130A
magscale 1 2
timestamp 1635355367
<< nwell >>
rect 91556 72130 92414 73734
rect 91554 71576 92414 72130
rect 91550 71320 92414 71576
rect 91550 71192 92412 71320
<< nmos >>
rect 91266 73478 91396 73514
rect 91108 73200 91396 73236
rect 90818 72784 91076 72820
rect 91294 72784 91394 72820
rect 90818 72512 91076 72548
rect 91294 72512 91394 72548
rect 90818 72240 91076 72276
rect 91294 72240 91394 72276
rect 90818 71968 91076 72004
rect 91292 71968 91392 72004
rect 90818 71696 91076 71732
rect 91292 71696 91392 71732
rect 90876 71366 91078 71402
<< pmos >>
rect 91610 73478 91868 73514
rect 91610 73200 92186 73236
rect 91610 72784 91710 72820
rect 91922 72786 92182 72822
rect 91610 72512 91710 72548
rect 91922 72514 92182 72550
rect 91610 72240 91710 72276
rect 91922 72242 92182 72278
rect 91608 71968 91708 72004
rect 91922 71970 92182 72006
rect 91608 71696 91708 71732
rect 91922 71698 92182 71734
rect 91922 71364 92124 71400
<< ndiff >>
rect 91266 73586 91396 73604
rect 91266 73550 91326 73586
rect 91362 73550 91396 73586
rect 91266 73514 91396 73550
rect 91266 73442 91396 73478
rect 91266 73406 91326 73442
rect 91362 73406 91396 73442
rect 91266 73388 91396 73406
rect 91108 73308 91396 73326
rect 91108 73272 91132 73308
rect 91166 73272 91206 73308
rect 91240 73272 91274 73308
rect 91308 73272 91344 73308
rect 91380 73272 91396 73308
rect 91108 73236 91396 73272
rect 91108 73164 91396 73200
rect 91108 73128 91132 73164
rect 91166 73128 91206 73164
rect 91240 73128 91274 73164
rect 91308 73128 91342 73164
rect 91378 73128 91396 73164
rect 91108 73110 91396 73128
rect 90818 72892 91076 72910
rect 90818 72856 90848 72892
rect 90882 72856 90922 72892
rect 90956 72856 91002 72892
rect 91036 72856 91076 72892
rect 91294 72892 91394 72910
rect 91294 72856 91326 72892
rect 91362 72856 91394 72892
rect 90818 72820 91076 72856
rect 91294 72820 91394 72856
rect 90818 72750 91076 72784
rect 90818 72748 91002 72750
rect 90818 72712 90848 72748
rect 90884 72712 90924 72748
rect 90960 72714 91002 72748
rect 91036 72714 91076 72750
rect 90960 72712 91076 72714
rect 90818 72694 91076 72712
rect 91294 72748 91394 72784
rect 91294 72712 91326 72748
rect 91362 72712 91394 72748
rect 91294 72694 91394 72712
rect 90818 72620 91076 72638
rect 90818 72584 90848 72620
rect 90882 72584 90922 72620
rect 90956 72584 91002 72620
rect 91036 72584 91076 72620
rect 91294 72620 91394 72638
rect 91294 72584 91326 72620
rect 91362 72584 91394 72620
rect 90818 72548 91076 72584
rect 91294 72548 91394 72584
rect 90818 72478 91076 72512
rect 90818 72476 91002 72478
rect 90818 72440 90848 72476
rect 90884 72440 90924 72476
rect 90960 72442 91002 72476
rect 91036 72442 91076 72478
rect 90960 72440 91076 72442
rect 90818 72422 91076 72440
rect 91294 72476 91394 72512
rect 91294 72440 91326 72476
rect 91362 72440 91394 72476
rect 91294 72422 91394 72440
rect 90818 72348 91076 72366
rect 90818 72312 90848 72348
rect 90882 72312 90922 72348
rect 90956 72312 91002 72348
rect 91036 72312 91076 72348
rect 91294 72348 91394 72366
rect 91294 72312 91326 72348
rect 91362 72312 91394 72348
rect 90818 72276 91076 72312
rect 91294 72276 91394 72312
rect 90818 72206 91076 72240
rect 90818 72204 91002 72206
rect 90818 72168 90848 72204
rect 90884 72168 90924 72204
rect 90960 72170 91002 72204
rect 91036 72170 91076 72206
rect 90960 72168 91076 72170
rect 90818 72150 91076 72168
rect 91294 72204 91394 72240
rect 91294 72168 91326 72204
rect 91362 72168 91394 72204
rect 91294 72150 91394 72168
rect 90818 72076 91076 72094
rect 90818 72040 90848 72076
rect 90882 72040 90922 72076
rect 90956 72040 91002 72076
rect 91036 72040 91076 72076
rect 91292 72076 91392 72094
rect 91292 72040 91324 72076
rect 91360 72040 91392 72076
rect 90818 72004 91076 72040
rect 91292 72004 91392 72040
rect 90818 71934 91076 71968
rect 90818 71932 91002 71934
rect 90818 71896 90848 71932
rect 90884 71896 90924 71932
rect 90960 71898 91002 71932
rect 91036 71898 91076 71934
rect 90960 71896 91076 71898
rect 90818 71878 91076 71896
rect 91292 71932 91392 71968
rect 91292 71896 91324 71932
rect 91360 71896 91392 71932
rect 91292 71878 91392 71896
rect 90818 71804 91076 71822
rect 90818 71768 90848 71804
rect 90882 71768 90922 71804
rect 90956 71768 91002 71804
rect 91036 71768 91076 71804
rect 91292 71804 91392 71822
rect 91292 71768 91324 71804
rect 91360 71768 91392 71804
rect 90818 71732 91076 71768
rect 91292 71732 91392 71768
rect 90818 71662 91076 71696
rect 90818 71660 91002 71662
rect 90818 71624 90848 71660
rect 90884 71624 90924 71660
rect 90960 71626 91002 71660
rect 91036 71626 91076 71662
rect 90960 71624 91076 71626
rect 90818 71606 91076 71624
rect 91292 71660 91392 71696
rect 91292 71624 91324 71660
rect 91360 71624 91392 71660
rect 91292 71606 91392 71624
rect 90876 71474 91078 71492
rect 90876 71438 90918 71474
rect 90952 71438 91002 71474
rect 91036 71438 91078 71474
rect 90876 71402 91078 71438
rect 90876 71330 91078 71366
rect 90876 71294 90920 71330
rect 90956 71294 91002 71330
rect 91038 71294 91078 71330
rect 90876 71276 91078 71294
<< pdiff >>
rect 91610 73586 91868 73604
rect 91610 73550 91642 73586
rect 91678 73550 91714 73586
rect 91750 73550 91784 73586
rect 91820 73550 91868 73586
rect 91610 73514 91868 73550
rect 91610 73442 91868 73478
rect 91610 73406 91642 73442
rect 91678 73406 91712 73442
rect 91748 73406 91782 73442
rect 91818 73406 91868 73442
rect 91610 73388 91868 73406
rect 91610 73310 92186 73326
rect 91610 73308 91712 73310
rect 91610 73272 91642 73308
rect 91678 73274 91712 73308
rect 91748 73274 91782 73310
rect 91818 73274 91852 73310
rect 91888 73274 91922 73310
rect 91958 73274 91992 73310
rect 92028 73274 92062 73310
rect 92098 73274 92132 73310
rect 92168 73274 92186 73310
rect 91678 73272 92186 73274
rect 91610 73236 92186 73272
rect 91610 73164 92186 73200
rect 91610 73128 91642 73164
rect 91678 73128 91712 73164
rect 91748 73128 91782 73164
rect 91818 73128 91852 73164
rect 91888 73128 91922 73164
rect 91958 73128 91992 73164
rect 92028 73128 92062 73164
rect 92098 73128 92132 73164
rect 92168 73128 92186 73164
rect 91610 73110 92186 73128
rect 91610 72892 91710 72910
rect 91610 72856 91642 72892
rect 91678 72856 91710 72892
rect 91922 72894 92182 72912
rect 91922 72858 91964 72894
rect 91998 72858 92044 72894
rect 92078 72858 92118 72894
rect 92152 72858 92182 72894
rect 91610 72820 91710 72856
rect 91922 72822 92182 72858
rect 91610 72748 91710 72784
rect 91610 72712 91642 72748
rect 91678 72712 91710 72748
rect 91610 72694 91710 72712
rect 91922 72752 92182 72786
rect 91922 72716 91964 72752
rect 91998 72750 92182 72752
rect 91998 72716 92040 72750
rect 91922 72714 92040 72716
rect 92076 72714 92116 72750
rect 92152 72714 92182 72750
rect 91922 72696 92182 72714
rect 91610 72620 91710 72638
rect 91610 72584 91642 72620
rect 91678 72584 91710 72620
rect 91922 72622 92182 72640
rect 91922 72586 91964 72622
rect 91998 72586 92044 72622
rect 92078 72586 92118 72622
rect 92152 72586 92182 72622
rect 91610 72548 91710 72584
rect 91922 72550 92182 72586
rect 91610 72476 91710 72512
rect 91610 72440 91642 72476
rect 91678 72440 91710 72476
rect 91610 72422 91710 72440
rect 91922 72480 92182 72514
rect 91922 72444 91964 72480
rect 91998 72478 92182 72480
rect 91998 72444 92040 72478
rect 91922 72442 92040 72444
rect 92076 72442 92116 72478
rect 92152 72442 92182 72478
rect 91922 72424 92182 72442
rect 91610 72348 91710 72366
rect 91610 72312 91642 72348
rect 91678 72312 91710 72348
rect 91922 72350 92182 72368
rect 91922 72314 91964 72350
rect 91998 72314 92044 72350
rect 92078 72314 92118 72350
rect 92152 72314 92182 72350
rect 91610 72276 91710 72312
rect 91922 72278 92182 72314
rect 91610 72204 91710 72240
rect 91610 72168 91642 72204
rect 91678 72168 91710 72204
rect 91610 72150 91710 72168
rect 91922 72208 92182 72242
rect 91922 72172 91964 72208
rect 91998 72206 92182 72208
rect 91998 72172 92040 72206
rect 91922 72170 92040 72172
rect 92076 72170 92116 72206
rect 92152 72170 92182 72206
rect 91922 72152 92182 72170
rect 91608 72076 91708 72094
rect 91608 72040 91640 72076
rect 91676 72040 91708 72076
rect 91922 72078 92182 72096
rect 91922 72042 91964 72078
rect 91998 72042 92044 72078
rect 92078 72042 92118 72078
rect 92152 72042 92182 72078
rect 91608 72004 91708 72040
rect 91922 72006 92182 72042
rect 91608 71932 91708 71968
rect 91608 71896 91640 71932
rect 91676 71896 91708 71932
rect 91608 71878 91708 71896
rect 91922 71936 92182 71970
rect 91922 71900 91964 71936
rect 91998 71934 92182 71936
rect 91998 71900 92040 71934
rect 91922 71898 92040 71900
rect 92076 71898 92116 71934
rect 92152 71898 92182 71934
rect 91922 71880 92182 71898
rect 91608 71804 91708 71822
rect 91608 71768 91640 71804
rect 91676 71768 91708 71804
rect 91922 71806 92182 71824
rect 91922 71770 91964 71806
rect 91998 71770 92044 71806
rect 92078 71770 92118 71806
rect 92152 71770 92182 71806
rect 91608 71732 91708 71768
rect 91922 71734 92182 71770
rect 91608 71660 91708 71696
rect 91608 71624 91640 71660
rect 91676 71624 91708 71660
rect 91608 71606 91708 71624
rect 91922 71664 92182 71698
rect 91922 71628 91964 71664
rect 91998 71662 92182 71664
rect 91998 71628 92040 71662
rect 91922 71626 92040 71628
rect 92076 71626 92116 71662
rect 92152 71626 92182 71662
rect 91922 71608 92182 71626
rect 91922 71474 92124 71490
rect 91922 71472 92024 71474
rect 91922 71436 91954 71472
rect 91990 71438 92024 71472
rect 92060 71438 92124 71474
rect 91990 71436 92124 71438
rect 91922 71400 92124 71436
rect 91922 71328 92124 71364
rect 91922 71292 91964 71328
rect 92000 71292 92046 71328
rect 92082 71292 92124 71328
rect 91922 71274 92124 71292
<< ndiffc >>
rect 91326 73550 91362 73586
rect 91326 73406 91362 73442
rect 91132 73272 91166 73308
rect 91206 73272 91240 73308
rect 91274 73272 91308 73308
rect 91344 73272 91380 73308
rect 91132 73128 91166 73164
rect 91206 73128 91240 73164
rect 91274 73128 91308 73164
rect 91342 73128 91378 73164
rect 90848 72856 90882 72892
rect 90922 72856 90956 72892
rect 91002 72856 91036 72892
rect 91326 72856 91362 72892
rect 90848 72712 90884 72748
rect 90924 72712 90960 72748
rect 91002 72714 91036 72750
rect 91326 72712 91362 72748
rect 90848 72584 90882 72620
rect 90922 72584 90956 72620
rect 91002 72584 91036 72620
rect 91326 72584 91362 72620
rect 90848 72440 90884 72476
rect 90924 72440 90960 72476
rect 91002 72442 91036 72478
rect 91326 72440 91362 72476
rect 90848 72312 90882 72348
rect 90922 72312 90956 72348
rect 91002 72312 91036 72348
rect 91326 72312 91362 72348
rect 90848 72168 90884 72204
rect 90924 72168 90960 72204
rect 91002 72170 91036 72206
rect 91326 72168 91362 72204
rect 90848 72040 90882 72076
rect 90922 72040 90956 72076
rect 91002 72040 91036 72076
rect 91324 72040 91360 72076
rect 90848 71896 90884 71932
rect 90924 71896 90960 71932
rect 91002 71898 91036 71934
rect 91324 71896 91360 71932
rect 90848 71768 90882 71804
rect 90922 71768 90956 71804
rect 91002 71768 91036 71804
rect 91324 71768 91360 71804
rect 90848 71624 90884 71660
rect 90924 71624 90960 71660
rect 91002 71626 91036 71662
rect 91324 71624 91360 71660
rect 90918 71438 90952 71474
rect 91002 71438 91036 71474
rect 90920 71294 90956 71330
rect 91002 71294 91038 71330
<< pdiffc >>
rect 91642 73550 91678 73586
rect 91714 73550 91750 73586
rect 91784 73550 91820 73586
rect 91642 73406 91678 73442
rect 91712 73406 91748 73442
rect 91782 73406 91818 73442
rect 91642 73272 91678 73308
rect 91712 73274 91748 73310
rect 91782 73274 91818 73310
rect 91852 73274 91888 73310
rect 91922 73274 91958 73310
rect 91992 73274 92028 73310
rect 92062 73274 92098 73310
rect 92132 73274 92168 73310
rect 91642 73128 91678 73164
rect 91712 73128 91748 73164
rect 91782 73128 91818 73164
rect 91852 73128 91888 73164
rect 91922 73128 91958 73164
rect 91992 73128 92028 73164
rect 92062 73128 92098 73164
rect 92132 73128 92168 73164
rect 91642 72856 91678 72892
rect 91964 72858 91998 72894
rect 92044 72858 92078 72894
rect 92118 72858 92152 72894
rect 91642 72712 91678 72748
rect 91964 72716 91998 72752
rect 92040 72714 92076 72750
rect 92116 72714 92152 72750
rect 91642 72584 91678 72620
rect 91964 72586 91998 72622
rect 92044 72586 92078 72622
rect 92118 72586 92152 72622
rect 91642 72440 91678 72476
rect 91964 72444 91998 72480
rect 92040 72442 92076 72478
rect 92116 72442 92152 72478
rect 91642 72312 91678 72348
rect 91964 72314 91998 72350
rect 92044 72314 92078 72350
rect 92118 72314 92152 72350
rect 91642 72168 91678 72204
rect 91964 72172 91998 72208
rect 92040 72170 92076 72206
rect 92116 72170 92152 72206
rect 91640 72040 91676 72076
rect 91964 72042 91998 72078
rect 92044 72042 92078 72078
rect 92118 72042 92152 72078
rect 91640 71896 91676 71932
rect 91964 71900 91998 71936
rect 92040 71898 92076 71934
rect 92116 71898 92152 71934
rect 91640 71768 91676 71804
rect 91964 71770 91998 71806
rect 92044 71770 92078 71806
rect 92118 71770 92152 71806
rect 91640 71624 91676 71660
rect 91964 71628 91998 71664
rect 92040 71626 92076 71662
rect 92116 71626 92152 71662
rect 91954 71436 91990 71472
rect 92024 71438 92060 71474
rect 91964 71292 92000 71328
rect 92046 71292 92082 71328
<< psubdiff >>
rect 90678 73322 90714 73346
rect 90678 73262 90714 73286
rect 90678 73046 90714 73070
rect 90678 72986 90714 73010
rect 90678 72704 90714 72728
rect 90678 72644 90714 72668
rect 90678 72430 90714 72454
rect 90678 72370 90714 72394
rect 90678 72158 90714 72182
rect 90678 72098 90714 72122
rect 90678 71888 90714 71912
rect 90678 71828 90714 71852
rect 90678 71566 90714 71590
rect 90678 71506 90714 71530
<< nsubdiff >>
rect 92284 73308 92320 73332
rect 92284 73248 92320 73272
rect 92284 73050 92320 73074
rect 92284 72990 92320 73014
rect 92284 72742 92320 72766
rect 92284 72682 92320 72706
rect 92284 72472 92320 72496
rect 92284 72412 92320 72436
rect 92284 72214 92320 72238
rect 92284 72154 92320 72178
rect 92276 71938 92326 71972
rect 92276 71902 92286 71938
rect 92322 71902 92326 71938
rect 92276 71874 92326 71902
rect 92286 71586 92322 71610
rect 92286 71526 92322 71550
<< psubdiffcont >>
rect 90678 73286 90714 73322
rect 90678 73010 90714 73046
rect 90678 72668 90714 72704
rect 90678 72394 90714 72430
rect 90678 72122 90714 72158
rect 90678 71852 90714 71888
rect 90678 71530 90714 71566
<< nsubdiffcont >>
rect 92284 73272 92320 73308
rect 92284 73014 92320 73050
rect 92284 72706 92320 72742
rect 92284 72436 92320 72472
rect 92284 72178 92320 72214
rect 92286 71902 92322 71938
rect 92286 71550 92322 71586
<< poly >>
rect 91240 73478 91266 73514
rect 91396 73490 91610 73514
rect 91396 73478 91490 73490
rect 91474 73454 91490 73478
rect 91526 73478 91610 73490
rect 91868 73478 91894 73514
rect 91526 73454 91542 73478
rect 91474 73440 91542 73454
rect 91486 73430 91530 73440
rect 91082 73200 91108 73236
rect 91396 73212 91610 73236
rect 91396 73200 91490 73212
rect 91474 73176 91490 73200
rect 91526 73200 91610 73212
rect 92186 73200 92212 73236
rect 91526 73176 91542 73200
rect 91474 73162 91542 73176
rect 91486 73152 91530 73162
rect 91122 72856 91166 72866
rect 91110 72842 91178 72856
rect 91110 72820 91126 72842
rect 90792 72784 90818 72820
rect 91076 72806 91126 72820
rect 91162 72806 91178 72842
rect 91834 72858 91878 72868
rect 91822 72844 91890 72858
rect 91076 72784 91178 72806
rect 91258 72784 91294 72820
rect 91394 72796 91610 72820
rect 91394 72784 91490 72796
rect 91474 72760 91490 72784
rect 91526 72784 91610 72796
rect 91710 72784 91746 72820
rect 91822 72808 91838 72844
rect 91874 72822 91890 72844
rect 91874 72808 91922 72822
rect 91822 72786 91922 72808
rect 92182 72786 92208 72822
rect 91526 72760 91542 72784
rect 91474 72746 91542 72760
rect 91486 72736 91530 72746
rect 91122 72584 91166 72594
rect 91110 72570 91178 72584
rect 91110 72548 91126 72570
rect 90792 72512 90818 72548
rect 91076 72534 91126 72548
rect 91162 72534 91178 72570
rect 91834 72586 91878 72596
rect 91822 72572 91890 72586
rect 91076 72512 91178 72534
rect 91258 72512 91294 72548
rect 91394 72524 91610 72548
rect 91394 72512 91490 72524
rect 91474 72488 91490 72512
rect 91526 72512 91610 72524
rect 91710 72512 91746 72548
rect 91822 72536 91838 72572
rect 91874 72550 91890 72572
rect 91874 72536 91922 72550
rect 91822 72514 91922 72536
rect 92182 72514 92208 72550
rect 91526 72488 91542 72512
rect 91474 72474 91542 72488
rect 91486 72464 91530 72474
rect 91122 72312 91166 72322
rect 91110 72298 91178 72312
rect 91110 72276 91126 72298
rect 90792 72240 90818 72276
rect 91076 72262 91126 72276
rect 91162 72262 91178 72298
rect 91834 72314 91878 72324
rect 91822 72300 91890 72314
rect 91076 72240 91178 72262
rect 91258 72240 91294 72276
rect 91394 72252 91610 72276
rect 91394 72240 91490 72252
rect 91474 72216 91490 72240
rect 91526 72240 91610 72252
rect 91710 72240 91746 72276
rect 91822 72264 91838 72300
rect 91874 72278 91890 72300
rect 91874 72264 91922 72278
rect 91822 72242 91922 72264
rect 92182 72242 92208 72278
rect 91526 72216 91542 72240
rect 91474 72202 91542 72216
rect 91486 72192 91530 72202
rect 91122 72040 91166 72050
rect 91110 72026 91178 72040
rect 91110 72004 91126 72026
rect 90792 71968 90818 72004
rect 91076 71990 91126 72004
rect 91162 71990 91178 72026
rect 91834 72042 91878 72052
rect 91822 72028 91890 72042
rect 91076 71968 91178 71990
rect 91256 71968 91292 72004
rect 91392 71980 91608 72004
rect 91392 71968 91488 71980
rect 91472 71944 91488 71968
rect 91524 71968 91608 71980
rect 91708 71968 91744 72004
rect 91822 71992 91838 72028
rect 91874 72006 91890 72028
rect 91874 71992 91922 72006
rect 91822 71970 91922 71992
rect 92182 71970 92208 72006
rect 91524 71944 91540 71968
rect 91472 71930 91540 71944
rect 91484 71920 91528 71930
rect 91122 71768 91166 71778
rect 91110 71754 91178 71768
rect 91110 71732 91126 71754
rect 90792 71696 90818 71732
rect 91076 71718 91126 71732
rect 91162 71718 91178 71754
rect 91834 71770 91878 71780
rect 91822 71756 91890 71770
rect 91076 71696 91178 71718
rect 91256 71696 91292 71732
rect 91392 71708 91608 71732
rect 91392 71696 91488 71708
rect 91472 71672 91488 71696
rect 91524 71696 91608 71708
rect 91708 71696 91744 71732
rect 91822 71720 91838 71756
rect 91874 71734 91890 71756
rect 91874 71720 91922 71734
rect 91822 71698 91922 71720
rect 92182 71698 92208 71734
rect 91524 71672 91540 71696
rect 91472 71658 91540 71672
rect 91484 71648 91528 71658
rect 91122 71438 91166 71448
rect 91110 71424 91178 71438
rect 91834 71436 91878 71446
rect 91110 71402 91126 71424
rect 90850 71366 90876 71402
rect 91078 71388 91126 71402
rect 91162 71388 91178 71424
rect 91078 71366 91178 71388
rect 91822 71422 91890 71436
rect 91822 71386 91838 71422
rect 91874 71400 91890 71422
rect 91874 71386 91922 71400
rect 91822 71364 91922 71386
rect 92124 71364 92150 71400
<< polycont >>
rect 91490 73454 91526 73490
rect 91490 73176 91526 73212
rect 91126 72806 91162 72842
rect 91490 72760 91526 72796
rect 91838 72808 91874 72844
rect 91126 72534 91162 72570
rect 91490 72488 91526 72524
rect 91838 72536 91874 72572
rect 91126 72262 91162 72298
rect 91490 72216 91526 72252
rect 91838 72264 91874 72300
rect 91126 71990 91162 72026
rect 91488 71944 91524 71980
rect 91838 71992 91874 72028
rect 91126 71718 91162 71754
rect 91488 71672 91524 71708
rect 91838 71720 91874 71756
rect 91126 71388 91162 71424
rect 91838 71386 91874 71422
<< locali >>
rect 91310 73590 91394 73602
rect 91490 73590 91526 73630
rect 91610 73590 91860 73602
rect 91310 73586 91860 73590
rect 91310 73550 91326 73586
rect 91362 73550 91642 73586
rect 91678 73550 91714 73586
rect 91750 73550 91784 73586
rect 91820 73550 91860 73586
rect 91310 73546 91860 73550
rect 91310 73534 91394 73546
rect 91610 73534 91860 73546
rect 90656 73456 90734 73500
rect 91474 73490 91542 73500
rect 91306 73456 91378 73458
rect 90656 73444 91378 73456
rect 91474 73454 91490 73490
rect 91526 73454 91542 73490
rect 92262 73458 92336 73472
rect 91474 73446 91542 73454
rect 90656 73408 90678 73444
rect 90714 73442 91378 73444
rect 90714 73408 91326 73442
rect 90656 73406 91326 73408
rect 91362 73406 91378 73442
rect 90656 73394 91378 73406
rect 90656 73322 90734 73394
rect 91306 73390 91378 73394
rect 90656 73286 90678 73322
rect 90714 73286 90734 73322
rect 90656 73180 90734 73286
rect 91124 73312 91394 73324
rect 91490 73312 91526 73446
rect 91622 73442 92336 73458
rect 91622 73406 91642 73442
rect 91678 73406 91712 73442
rect 91748 73406 91782 73442
rect 91818 73406 92282 73442
rect 92318 73406 92336 73442
rect 91622 73390 92336 73406
rect 91610 73320 91692 73324
rect 91610 73312 92184 73320
rect 91124 73310 92184 73312
rect 91124 73308 91712 73310
rect 91124 73272 91132 73308
rect 91166 73272 91206 73308
rect 91240 73272 91274 73308
rect 91308 73272 91344 73308
rect 91380 73272 91642 73308
rect 91678 73274 91712 73308
rect 91748 73274 91782 73310
rect 91818 73274 91852 73310
rect 91888 73274 91922 73310
rect 91958 73274 91992 73310
rect 92028 73274 92062 73310
rect 92098 73274 92132 73310
rect 92168 73274 92184 73310
rect 91678 73272 92184 73274
rect 91124 73268 92184 73272
rect 91124 73258 91394 73268
rect 91132 73256 91394 73258
rect 91610 73256 92184 73268
rect 92262 73308 92336 73390
rect 92262 73272 92284 73308
rect 92320 73272 92336 73308
rect 91474 73212 91542 73222
rect 90656 73164 91392 73180
rect 91474 73176 91490 73212
rect 91526 73176 91542 73212
rect 92262 73182 92336 73272
rect 92164 73180 92336 73182
rect 91474 73168 91542 73176
rect 90656 73158 91132 73164
rect 90656 73122 90678 73158
rect 90714 73128 91132 73158
rect 91166 73128 91206 73164
rect 91240 73128 91274 73164
rect 91308 73128 91342 73164
rect 91378 73128 91392 73164
rect 90714 73122 91392 73128
rect 90656 73114 91392 73122
rect 90656 73112 91378 73114
rect 90656 73046 90734 73112
rect 90656 73010 90678 73046
rect 90714 73010 90734 73046
rect 90656 72906 90734 73010
rect 91490 72964 91526 73168
rect 91622 73166 92336 73180
rect 91622 73164 92282 73166
rect 91622 73128 91642 73164
rect 91678 73128 91712 73164
rect 91748 73128 91782 73164
rect 91818 73128 91852 73164
rect 91888 73128 91922 73164
rect 91958 73128 91992 73164
rect 92028 73128 92062 73164
rect 92098 73128 92132 73164
rect 92168 73130 92282 73164
rect 92318 73130 92336 73166
rect 92168 73128 92336 73130
rect 91622 73114 92336 73128
rect 91622 73112 92178 73114
rect 92262 73050 92336 73114
rect 92262 73014 92284 73050
rect 92320 73014 92336 73050
rect 90818 72906 91062 72908
rect 90656 72892 91062 72906
rect 90656 72890 90848 72892
rect 90656 72854 90678 72890
rect 90714 72856 90848 72890
rect 90882 72856 90922 72892
rect 90956 72856 91002 72892
rect 91036 72856 91062 72892
rect 90714 72854 91062 72856
rect 90656 72842 91062 72854
rect 91126 72850 91162 72884
rect 91310 72896 91394 72908
rect 91490 72896 91526 72922
rect 91610 72896 91692 72908
rect 91310 72892 91692 72896
rect 91310 72856 91326 72892
rect 91362 72856 91642 72892
rect 91678 72856 91692 72892
rect 91310 72852 91692 72856
rect 92262 72912 92336 73014
rect 92178 72910 92336 72912
rect 91838 72852 91874 72886
rect 91938 72906 92336 72910
rect 91938 72896 92338 72906
rect 91938 72894 92282 72896
rect 91938 72858 91964 72894
rect 91998 72858 92044 72894
rect 92078 72858 92118 72894
rect 92152 72860 92282 72894
rect 92318 72860 92338 72896
rect 92152 72858 92338 72860
rect 90656 72704 90734 72842
rect 90818 72840 91062 72842
rect 91110 72842 91178 72850
rect 91110 72806 91126 72842
rect 91162 72806 91178 72842
rect 91310 72840 91394 72852
rect 91610 72840 91692 72852
rect 91822 72844 91890 72852
rect 91822 72808 91838 72844
rect 91874 72808 91890 72844
rect 91938 72844 92338 72858
rect 91938 72842 92182 72844
rect 91110 72796 91178 72806
rect 91474 72796 91542 72806
rect 91822 72798 91890 72808
rect 90656 72668 90678 72704
rect 90714 72668 90734 72704
rect 90818 72754 91076 72766
rect 90818 72752 91078 72754
rect 91306 72752 91378 72764
rect 91474 72760 91490 72796
rect 91526 72760 91542 72796
rect 91474 72752 91542 72760
rect 91622 72754 91694 72764
rect 91924 72756 92182 72768
rect 91922 72754 92182 72756
rect 91622 72752 92182 72754
rect 90818 72750 91378 72752
rect 90818 72748 91002 72750
rect 90818 72712 90848 72748
rect 90884 72712 90924 72748
rect 90960 72714 91002 72748
rect 91036 72748 91378 72750
rect 91036 72714 91326 72748
rect 90960 72712 91326 72714
rect 91362 72712 91378 72748
rect 90818 72706 91378 72712
rect 90818 72696 91076 72706
rect 91306 72696 91378 72706
rect 90656 72634 90734 72668
rect 90818 72634 91062 72636
rect 90656 72620 91062 72634
rect 90656 72584 90848 72620
rect 90882 72584 90922 72620
rect 90956 72584 91002 72620
rect 91036 72584 91062 72620
rect 90656 72570 91062 72584
rect 91126 72578 91162 72612
rect 91310 72624 91394 72636
rect 91490 72624 91526 72752
rect 91622 72748 91964 72752
rect 91622 72712 91642 72748
rect 91678 72716 91964 72748
rect 91998 72750 92182 72752
rect 91998 72716 92040 72750
rect 91678 72714 92040 72716
rect 92076 72714 92116 72750
rect 92152 72714 92182 72750
rect 91678 72712 92182 72714
rect 91622 72708 92182 72712
rect 91622 72696 91694 72708
rect 91924 72698 92182 72708
rect 92262 72742 92338 72844
rect 92262 72706 92284 72742
rect 92320 72706 92338 72742
rect 91610 72624 91692 72636
rect 91310 72620 91692 72624
rect 91310 72584 91326 72620
rect 91362 72584 91642 72620
rect 91678 72584 91692 72620
rect 91310 72580 91692 72584
rect 92262 72640 92338 72706
rect 92180 72638 92338 72640
rect 91838 72580 91874 72614
rect 91938 72622 92338 72638
rect 91938 72586 91964 72622
rect 91998 72586 92044 72622
rect 92078 72586 92118 72622
rect 92152 72586 92284 72622
rect 92320 72586 92338 72622
rect 90656 72534 90678 72570
rect 90714 72534 90734 72570
rect 90818 72568 91062 72570
rect 91110 72570 91178 72578
rect 90656 72430 90734 72534
rect 91110 72534 91126 72570
rect 91162 72534 91178 72570
rect 91310 72568 91394 72580
rect 91610 72568 91692 72580
rect 91822 72572 91890 72580
rect 91822 72536 91838 72572
rect 91874 72536 91890 72572
rect 91938 72572 92338 72586
rect 91938 72570 92182 72572
rect 91110 72524 91178 72534
rect 91474 72524 91542 72534
rect 91822 72526 91890 72536
rect 90656 72394 90678 72430
rect 90714 72394 90734 72430
rect 90818 72482 91076 72494
rect 90818 72480 91078 72482
rect 91306 72480 91378 72492
rect 91474 72488 91490 72524
rect 91526 72488 91542 72524
rect 91474 72480 91542 72488
rect 91622 72482 91694 72492
rect 91924 72484 92182 72496
rect 91922 72482 92182 72484
rect 91622 72480 92182 72482
rect 90818 72478 91378 72480
rect 90818 72476 91002 72478
rect 90818 72440 90848 72476
rect 90884 72440 90924 72476
rect 90960 72442 91002 72476
rect 91036 72476 91378 72478
rect 91036 72442 91326 72476
rect 90960 72440 91326 72442
rect 91362 72440 91378 72476
rect 90818 72434 91378 72440
rect 90818 72424 91076 72434
rect 91306 72424 91378 72434
rect 90656 72364 90734 72394
rect 90656 72348 91062 72364
rect 90656 72312 90848 72348
rect 90882 72312 90922 72348
rect 90956 72312 91002 72348
rect 91036 72312 91062 72348
rect 90656 72300 91062 72312
rect 91126 72306 91162 72340
rect 91310 72352 91394 72364
rect 91490 72352 91526 72480
rect 91622 72476 91964 72480
rect 91622 72440 91642 72476
rect 91678 72444 91964 72476
rect 91998 72478 92182 72480
rect 91998 72444 92040 72478
rect 91678 72442 92040 72444
rect 92076 72442 92116 72478
rect 92152 72442 92182 72478
rect 91678 72440 92182 72442
rect 91622 72436 92182 72440
rect 91622 72424 91694 72436
rect 91924 72426 92182 72436
rect 92262 72472 92338 72572
rect 92262 72436 92284 72472
rect 92320 72436 92338 72472
rect 91610 72352 91692 72364
rect 91310 72348 91692 72352
rect 91310 72312 91326 72348
rect 91362 72312 91642 72348
rect 91678 72312 91692 72348
rect 91310 72308 91692 72312
rect 92262 72366 92338 72436
rect 91838 72308 91874 72342
rect 91938 72350 92338 72366
rect 91938 72314 91964 72350
rect 91998 72314 92044 72350
rect 92078 72314 92118 72350
rect 92152 72314 92286 72350
rect 92322 72314 92338 72350
rect 90656 72294 90734 72300
rect 90818 72296 91062 72300
rect 91110 72298 91178 72306
rect 90656 72258 90678 72294
rect 90714 72258 90734 72294
rect 90656 72158 90734 72258
rect 91110 72262 91126 72298
rect 91162 72262 91178 72298
rect 91310 72296 91394 72308
rect 91610 72296 91692 72308
rect 91822 72300 91890 72308
rect 91822 72264 91838 72300
rect 91874 72264 91890 72300
rect 91938 72298 92338 72314
rect 91110 72252 91178 72262
rect 91474 72252 91542 72262
rect 91822 72254 91890 72264
rect 90656 72122 90678 72158
rect 90714 72122 90734 72158
rect 90818 72210 91076 72222
rect 90818 72208 91078 72210
rect 91306 72208 91378 72220
rect 91474 72216 91490 72252
rect 91526 72216 91542 72252
rect 91474 72208 91542 72216
rect 91622 72210 91694 72220
rect 91924 72212 92182 72224
rect 91922 72210 92182 72212
rect 91622 72208 92182 72210
rect 90818 72206 91378 72208
rect 90818 72204 91002 72206
rect 90818 72168 90848 72204
rect 90884 72168 90924 72204
rect 90960 72170 91002 72204
rect 91036 72204 91378 72206
rect 91036 72170 91326 72204
rect 90960 72168 91326 72170
rect 91362 72168 91378 72204
rect 90818 72162 91378 72168
rect 90818 72152 91076 72162
rect 91306 72152 91378 72162
rect 91490 72160 91526 72208
rect 90656 72090 90734 72122
rect 91488 72132 91526 72160
rect 91622 72204 91964 72208
rect 91622 72168 91642 72204
rect 91678 72172 91964 72204
rect 91998 72206 92182 72208
rect 91998 72172 92040 72206
rect 91678 72170 92040 72172
rect 92076 72170 92116 72206
rect 92152 72170 92182 72206
rect 91678 72168 92182 72170
rect 91622 72164 92182 72168
rect 91622 72152 91694 72164
rect 91924 72154 92182 72164
rect 92262 72214 92338 72298
rect 92262 72178 92284 72214
rect 92320 72178 92338 72214
rect 90818 72090 91062 72092
rect 90656 72076 91062 72090
rect 90656 72040 90848 72076
rect 90882 72040 90922 72076
rect 90956 72040 91002 72076
rect 91036 72040 91062 72076
rect 90656 72026 91062 72040
rect 91126 72034 91162 72068
rect 91308 72080 91392 72092
rect 91488 72080 91524 72132
rect 91608 72080 91690 72092
rect 91308 72076 91690 72080
rect 91308 72040 91324 72076
rect 91360 72040 91640 72076
rect 91676 72040 91690 72076
rect 91308 72036 91690 72040
rect 92262 72094 92338 72178
rect 91838 72036 91874 72070
rect 91938 72080 92338 72094
rect 91938 72078 92286 72080
rect 91938 72042 91964 72078
rect 91998 72042 92044 72078
rect 92078 72042 92118 72078
rect 92152 72044 92286 72078
rect 92322 72044 92338 72080
rect 92152 72042 92338 72044
rect 90656 72022 90734 72026
rect 90818 72024 91062 72026
rect 91110 72026 91178 72034
rect 90656 71986 90678 72022
rect 90714 71986 90734 72022
rect 90656 71888 90734 71986
rect 91110 71990 91126 72026
rect 91162 71990 91178 72026
rect 91308 72024 91392 72036
rect 91608 72024 91690 72036
rect 91822 72028 91890 72036
rect 91822 71992 91838 72028
rect 91874 71992 91890 72028
rect 91938 72026 92338 72042
rect 91110 71980 91178 71990
rect 91472 71980 91540 71990
rect 91822 71982 91890 71992
rect 90656 71852 90678 71888
rect 90714 71852 90734 71888
rect 90818 71938 91076 71950
rect 90818 71936 91078 71938
rect 91304 71936 91376 71948
rect 91472 71944 91488 71980
rect 91524 71944 91540 71980
rect 91472 71936 91540 71944
rect 91620 71938 91692 71948
rect 91924 71940 92182 71952
rect 91922 71938 92182 71940
rect 91620 71936 92182 71938
rect 90818 71934 91376 71936
rect 90818 71932 91002 71934
rect 90818 71896 90848 71932
rect 90884 71896 90924 71932
rect 90960 71898 91002 71932
rect 91036 71932 91376 71934
rect 91036 71898 91324 71932
rect 90960 71896 91324 71898
rect 91360 71896 91376 71932
rect 90818 71890 91376 71896
rect 90818 71880 91076 71890
rect 91304 71880 91376 71890
rect 90656 71818 90734 71852
rect 90818 71818 91062 71820
rect 90656 71804 91062 71818
rect 90656 71768 90848 71804
rect 90882 71768 90922 71804
rect 90956 71768 91002 71804
rect 91036 71768 91062 71804
rect 90656 71754 91062 71768
rect 91126 71762 91162 71796
rect 91308 71808 91392 71820
rect 91488 71808 91524 71936
rect 91620 71932 91964 71936
rect 91620 71896 91640 71932
rect 91676 71900 91964 71932
rect 91998 71934 92182 71936
rect 91998 71900 92040 71934
rect 91676 71898 92040 71900
rect 92076 71898 92116 71934
rect 92152 71898 92182 71934
rect 91676 71896 92182 71898
rect 91620 71892 92182 71896
rect 91620 71880 91692 71892
rect 91924 71882 92182 71892
rect 92262 71938 92338 72026
rect 92262 71902 92286 71938
rect 92322 71902 92338 71938
rect 91608 71808 91690 71820
rect 91308 71804 91690 71808
rect 91308 71768 91324 71804
rect 91360 71768 91640 71804
rect 91676 71768 91690 71804
rect 91308 71764 91690 71768
rect 92262 71824 92338 71902
rect 92182 71822 92338 71824
rect 91838 71764 91874 71798
rect 91938 71808 92338 71822
rect 91938 71806 92286 71808
rect 91938 71770 91964 71806
rect 91998 71770 92044 71806
rect 92078 71770 92118 71806
rect 92152 71772 92286 71806
rect 92322 71772 92338 71808
rect 92152 71770 92338 71772
rect 90656 71710 90734 71754
rect 90818 71752 91062 71754
rect 91110 71754 91178 71762
rect 90656 71674 90678 71710
rect 90714 71674 90734 71710
rect 91110 71718 91126 71754
rect 91162 71718 91178 71754
rect 91308 71752 91392 71764
rect 91608 71752 91690 71764
rect 91822 71756 91890 71764
rect 91822 71720 91838 71756
rect 91874 71720 91890 71756
rect 91938 71756 92338 71770
rect 91938 71754 92182 71756
rect 92262 71754 92338 71756
rect 91110 71708 91178 71718
rect 91472 71708 91540 71718
rect 91822 71710 91890 71720
rect 90656 71566 90734 71674
rect 90818 71666 91076 71678
rect 90818 71664 91078 71666
rect 91304 71664 91376 71676
rect 91472 71672 91488 71708
rect 91524 71672 91540 71708
rect 91472 71664 91540 71672
rect 91620 71666 91692 71676
rect 91924 71668 92182 71680
rect 91922 71666 92182 71668
rect 91620 71664 92182 71666
rect 90818 71662 91376 71664
rect 90818 71660 91002 71662
rect 90818 71624 90848 71660
rect 90884 71624 90924 71660
rect 90960 71626 91002 71660
rect 91036 71660 91376 71662
rect 91036 71626 91324 71660
rect 90960 71624 91324 71626
rect 91360 71624 91376 71660
rect 90818 71618 91376 71624
rect 90818 71608 91076 71618
rect 91304 71608 91376 71618
rect 91488 71630 91524 71664
rect 91620 71660 91964 71664
rect 91620 71624 91640 71660
rect 91676 71628 91964 71660
rect 91998 71662 92182 71664
rect 91998 71628 92040 71662
rect 91676 71626 92040 71628
rect 92076 71626 92116 71662
rect 92152 71626 92182 71662
rect 91676 71624 92182 71626
rect 91620 71620 92182 71624
rect 91620 71608 91692 71620
rect 91924 71610 92182 71620
rect 90656 71530 90678 71566
rect 90714 71530 90734 71566
rect 90656 71484 90734 71530
rect 92264 71586 92338 71754
rect 92264 71550 92286 71586
rect 92322 71550 92338 71586
rect 90876 71484 91058 71490
rect 90656 71474 91058 71484
rect 90656 71472 90918 71474
rect 90656 71436 90678 71472
rect 90714 71438 90918 71472
rect 90952 71438 91002 71474
rect 91036 71438 91058 71474
rect 90714 71436 91058 71438
rect 90656 71430 91058 71436
rect 91126 71432 91162 71466
rect 92264 71484 92338 71550
rect 90656 71370 90734 71430
rect 90876 71422 91058 71430
rect 91110 71424 91178 71432
rect 91838 71430 91874 71464
rect 91934 71474 92338 71484
rect 91934 71472 92024 71474
rect 91934 71436 91954 71472
rect 91990 71438 92024 71472
rect 92060 71468 92338 71474
rect 92060 71438 92286 71468
rect 91990 71436 92286 71438
rect 91934 71432 92286 71436
rect 92322 71432 92338 71468
rect 91110 71388 91126 71424
rect 91162 71388 91178 71424
rect 91110 71378 91178 71388
rect 91822 71422 91890 71430
rect 91822 71386 91838 71422
rect 91874 71386 91890 71422
rect 91934 71420 92338 71432
rect 91822 71376 91890 71386
rect 90876 71336 91058 71348
rect 91828 71340 91878 71376
rect 91926 71340 92106 71344
rect 91828 71336 92106 71340
rect 90876 71330 92106 71336
rect 90876 71294 90920 71330
rect 90956 71294 91002 71330
rect 91038 71328 92106 71330
rect 91038 71294 91964 71328
rect 90876 71292 91964 71294
rect 92000 71292 92046 71328
rect 92082 71292 92106 71328
rect 90876 71284 92106 71292
rect 90876 71278 91058 71284
rect 91828 71282 92106 71284
rect 91922 71276 92106 71282
rect 92264 71186 92338 71420
rect 92264 70996 92336 71186
rect 92266 70830 92336 70996
rect 92266 70792 92282 70830
rect 92320 70792 92336 70830
rect 92266 70782 92336 70792
<< viali >>
rect 91490 73630 91526 73666
rect 90678 73408 90714 73444
rect 92282 73406 92318 73442
rect 90678 73122 90714 73158
rect 92282 73130 92318 73166
rect 91490 72922 91526 72964
rect 90678 72854 90714 72890
rect 91126 72884 91162 72922
rect 91838 72886 91874 72924
rect 92282 72860 92318 72896
rect 91126 72612 91162 72650
rect 91838 72614 91874 72652
rect 92284 72586 92320 72622
rect 90678 72534 90714 72570
rect 91126 72340 91162 72378
rect 91838 72342 91874 72380
rect 92286 72314 92322 72350
rect 90678 72258 90714 72294
rect 91126 72068 91162 72106
rect 91838 72070 91874 72108
rect 92286 72044 92322 72080
rect 90678 71986 90714 72022
rect 91126 71796 91162 71834
rect 91838 71798 91874 71836
rect 92286 71772 92322 71808
rect 90678 71674 90714 71710
rect 91488 71588 91524 71630
rect 90678 71436 90714 71472
rect 91126 71466 91162 71504
rect 91838 71464 91874 71502
rect 92286 71432 92322 71468
rect 92282 70792 92320 70830
<< metal1 >>
rect 91474 73820 91544 73900
rect 91470 73810 91548 73820
rect 91470 73754 91482 73810
rect 91538 73754 91548 73810
rect 91470 73734 91548 73754
rect 91478 73666 91536 73734
rect 90660 73582 90730 73662
rect 91478 73630 91490 73666
rect 91526 73630 91536 73666
rect 91478 73600 91536 73630
rect 90656 73572 90734 73582
rect 90656 73516 90668 73572
rect 90724 73516 90734 73572
rect 90656 73500 90734 73516
rect 90654 73496 90734 73500
rect 90654 73444 90736 73496
rect 90654 73408 90678 73444
rect 90714 73408 90736 73444
rect 90654 73158 90736 73408
rect 90654 73122 90678 73158
rect 90714 73122 90736 73158
rect 90654 72890 90736 73122
rect 92266 73442 92338 73470
rect 92266 73406 92282 73442
rect 92318 73406 92338 73442
rect 92266 73166 92338 73406
rect 92266 73130 92282 73166
rect 92318 73130 92338 73166
rect 91478 72964 91536 72976
rect 90654 72854 90678 72890
rect 90714 72854 90736 72890
rect 90654 72570 90736 72854
rect 90654 72534 90678 72570
rect 90714 72534 90736 72570
rect 90654 72294 90736 72534
rect 90654 72258 90678 72294
rect 90714 72258 90736 72294
rect 90654 72022 90736 72258
rect 90654 71986 90678 72022
rect 90714 71986 90736 72022
rect 90654 71710 90736 71986
rect 90654 71674 90678 71710
rect 90714 71674 90736 71710
rect 90654 71472 90736 71674
rect 90654 71436 90678 71472
rect 90714 71436 90736 71472
rect 90654 71368 90736 71436
rect 91116 72922 91174 72936
rect 91116 72884 91126 72922
rect 91162 72884 91174 72922
rect 91116 72650 91174 72884
rect 91116 72612 91126 72650
rect 91162 72612 91174 72650
rect 91116 72378 91174 72612
rect 91116 72340 91126 72378
rect 91162 72340 91174 72378
rect 91116 72106 91174 72340
rect 91116 72068 91126 72106
rect 91162 72068 91174 72106
rect 91116 71834 91174 72068
rect 91116 71796 91126 71834
rect 91162 71796 91174 71834
rect 91116 71504 91174 71796
rect 91478 72922 91490 72964
rect 91526 72922 91536 72964
rect 91478 71630 91536 72922
rect 91478 71588 91488 71630
rect 91524 71588 91536 71630
rect 91478 71561 91536 71588
rect 91826 72924 91884 72938
rect 91826 72886 91838 72924
rect 91874 72886 91884 72924
rect 91826 72652 91884 72886
rect 91826 72614 91838 72652
rect 91874 72614 91884 72652
rect 91826 72380 91884 72614
rect 91826 72342 91838 72380
rect 91874 72342 91884 72380
rect 91826 72108 91884 72342
rect 91826 72070 91838 72108
rect 91874 72070 91884 72108
rect 91826 71836 91884 72070
rect 91826 71798 91838 71836
rect 91874 71798 91884 71836
rect 91116 71466 91126 71504
rect 91162 71466 91174 71504
rect 91116 71438 91174 71466
rect 91826 71502 91884 71798
rect 92266 72896 92338 73130
rect 92266 72860 92282 72896
rect 92318 72860 92338 72896
rect 92266 72622 92338 72860
rect 92266 72586 92284 72622
rect 92320 72586 92338 72622
rect 92266 72350 92338 72586
rect 92266 72314 92286 72350
rect 92322 72314 92338 72350
rect 92266 72080 92338 72314
rect 92266 72044 92286 72080
rect 92322 72044 92338 72080
rect 92266 71808 92338 72044
rect 92266 71772 92286 71808
rect 92322 71772 92338 71808
rect 92266 71748 92338 71772
rect 91826 71464 91838 71502
rect 91874 71464 91884 71502
rect 91116 71437 91226 71438
rect 91116 71367 91536 71437
rect 91116 71366 91226 71367
rect 91478 71105 91536 71367
rect 91826 71364 91884 71464
rect 92264 71468 92338 71748
rect 92264 71432 92286 71468
rect 92322 71432 92338 71468
rect 92264 71368 92338 71432
rect 91478 71025 91537 71105
rect 91471 70917 91549 71025
rect 91471 70861 91481 70917
rect 91537 70861 91549 70917
rect 91471 70851 91549 70861
rect 91475 70771 91545 70851
rect 92268 70830 92334 70846
rect 92268 70792 92282 70830
rect 92320 70792 92334 70830
rect 92268 70784 92334 70792
rect 92272 70736 92330 70784
rect 92260 70716 92338 70736
rect 92260 70660 92270 70716
rect 92326 70660 92338 70716
rect 92260 70650 92338 70660
rect 92264 70570 92334 70650
<< via1 >>
rect 91482 73754 91538 73810
rect 90668 73516 90724 73572
rect 91481 70861 91537 70917
rect 92270 70660 92326 70716
<< metal2 >>
rect 91474 73820 91544 73900
rect 91470 73810 91548 73820
rect 91470 73754 91482 73810
rect 91538 73754 91548 73810
rect 91470 73734 91548 73754
rect 90660 73582 90730 73662
rect 90656 73572 90734 73582
rect 90656 73516 90668 73572
rect 90724 73516 90734 73572
rect 90656 73496 90734 73516
rect 91471 70917 91549 70937
rect 91471 70861 91481 70917
rect 91537 70861 91549 70917
rect 91471 70851 91549 70861
rect 91475 70771 91545 70851
rect 92260 70716 92338 70736
rect 92260 70660 92270 70716
rect 92326 70660 92338 70716
rect 92260 70650 92338 70660
rect 92264 70570 92334 70650
<< via2 >>
rect 91482 73754 91538 73810
rect 90668 73516 90724 73572
rect 91481 70861 91537 70917
rect 92270 70660 92326 70716
<< metal3 >>
rect 66138 93042 66896 93112
rect -38198 92953 -37486 93024
rect 14114 92964 14954 93034
rect -37810 69255 -37739 92953
rect 14516 70580 14586 92964
rect 66538 73853 66608 93042
rect 111216 92928 111882 92998
rect 91474 75414 91544 75466
rect 111512 75414 111582 92928
rect 91474 75344 111610 75414
rect 66538 73783 90730 73853
rect 91474 73820 91544 75344
rect 111512 75311 111582 75344
rect 90660 73582 90730 73783
rect 91470 73810 91548 73820
rect 91470 73754 91482 73810
rect 91538 73754 91548 73810
rect 91470 73734 91548 73754
rect 90656 73572 90734 73582
rect 90656 73516 90668 73572
rect 90724 73516 90734 73572
rect 90656 73496 90734 73516
rect 91471 70917 91549 70937
rect 91471 70861 91481 70917
rect 91537 70861 91549 70917
rect 91471 70851 91549 70861
rect 91475 70580 91545 70851
rect 92260 70716 92338 70736
rect 92260 70660 92270 70716
rect 92326 70660 92338 70716
rect 92260 70650 92338 70660
rect 14516 70510 91545 70580
rect 92264 70585 92334 70650
rect 92264 69255 92335 70585
rect -37810 69184 92335 69255
<< labels >>
rlabel metal3 92299 70605 92299 70605 1 io_analog[9]
rlabel metal3 91509 70805 91509 70805 1 io_analog[8]
rlabel metal3 90697 73621 90697 73621 1 io_analog[7]
rlabel metal3 91509 73857 91509 73857 1 io_analog[6]
<< end >>
