magic
tech sky130A
magscale 1 2
timestamp 1633447108
<< nwell >>
rect 31556 32130 32414 33734
rect 31554 31576 32414 32130
rect 31550 31320 32414 31576
rect 31550 31192 32412 31320
<< nmos >>
rect 31266 33478 31396 33514
rect 31108 33200 31396 33236
rect 30818 32784 31076 32820
rect 31294 32784 31394 32820
rect 30818 32512 31076 32548
rect 31294 32512 31394 32548
rect 30818 32240 31076 32276
rect 31294 32240 31394 32276
rect 30818 31968 31076 32004
rect 31292 31968 31392 32004
rect 30818 31696 31076 31732
rect 31292 31696 31392 31732
rect 30876 31366 31078 31402
<< pmos >>
rect 31610 33478 31868 33514
rect 31610 33200 32186 33236
rect 31610 32784 31710 32820
rect 31922 32786 32182 32822
rect 31610 32512 31710 32548
rect 31922 32514 32182 32550
rect 31610 32240 31710 32276
rect 31922 32242 32182 32278
rect 31608 31968 31708 32004
rect 31922 31970 32182 32006
rect 31608 31696 31708 31732
rect 31922 31698 32182 31734
rect 31922 31364 32124 31400
<< ndiff >>
rect 31266 33586 31396 33604
rect 31266 33550 31326 33586
rect 31362 33550 31396 33586
rect 31266 33514 31396 33550
rect 31266 33442 31396 33478
rect 31266 33406 31326 33442
rect 31362 33406 31396 33442
rect 31266 33388 31396 33406
rect 31108 33308 31396 33326
rect 31108 33272 31132 33308
rect 31166 33272 31206 33308
rect 31240 33272 31274 33308
rect 31308 33272 31344 33308
rect 31380 33272 31396 33308
rect 31108 33236 31396 33272
rect 31108 33164 31396 33200
rect 31108 33128 31132 33164
rect 31166 33128 31206 33164
rect 31240 33128 31274 33164
rect 31308 33128 31342 33164
rect 31378 33128 31396 33164
rect 31108 33110 31396 33128
rect 30818 32892 31076 32910
rect 30818 32856 30848 32892
rect 30882 32856 30922 32892
rect 30956 32856 31002 32892
rect 31036 32856 31076 32892
rect 31294 32892 31394 32910
rect 31294 32856 31326 32892
rect 31362 32856 31394 32892
rect 30818 32820 31076 32856
rect 31294 32820 31394 32856
rect 30818 32750 31076 32784
rect 30818 32748 31002 32750
rect 30818 32712 30848 32748
rect 30884 32712 30924 32748
rect 30960 32714 31002 32748
rect 31036 32714 31076 32750
rect 30960 32712 31076 32714
rect 30818 32694 31076 32712
rect 31294 32748 31394 32784
rect 31294 32712 31326 32748
rect 31362 32712 31394 32748
rect 31294 32694 31394 32712
rect 30818 32620 31076 32638
rect 30818 32584 30848 32620
rect 30882 32584 30922 32620
rect 30956 32584 31002 32620
rect 31036 32584 31076 32620
rect 31294 32620 31394 32638
rect 31294 32584 31326 32620
rect 31362 32584 31394 32620
rect 30818 32548 31076 32584
rect 31294 32548 31394 32584
rect 30818 32478 31076 32512
rect 30818 32476 31002 32478
rect 30818 32440 30848 32476
rect 30884 32440 30924 32476
rect 30960 32442 31002 32476
rect 31036 32442 31076 32478
rect 30960 32440 31076 32442
rect 30818 32422 31076 32440
rect 31294 32476 31394 32512
rect 31294 32440 31326 32476
rect 31362 32440 31394 32476
rect 31294 32422 31394 32440
rect 30818 32348 31076 32366
rect 30818 32312 30848 32348
rect 30882 32312 30922 32348
rect 30956 32312 31002 32348
rect 31036 32312 31076 32348
rect 31294 32348 31394 32366
rect 31294 32312 31326 32348
rect 31362 32312 31394 32348
rect 30818 32276 31076 32312
rect 31294 32276 31394 32312
rect 30818 32206 31076 32240
rect 30818 32204 31002 32206
rect 30818 32168 30848 32204
rect 30884 32168 30924 32204
rect 30960 32170 31002 32204
rect 31036 32170 31076 32206
rect 30960 32168 31076 32170
rect 30818 32150 31076 32168
rect 31294 32204 31394 32240
rect 31294 32168 31326 32204
rect 31362 32168 31394 32204
rect 31294 32150 31394 32168
rect 30818 32076 31076 32094
rect 30818 32040 30848 32076
rect 30882 32040 30922 32076
rect 30956 32040 31002 32076
rect 31036 32040 31076 32076
rect 31292 32076 31392 32094
rect 31292 32040 31324 32076
rect 31360 32040 31392 32076
rect 30818 32004 31076 32040
rect 31292 32004 31392 32040
rect 30818 31934 31076 31968
rect 30818 31932 31002 31934
rect 30818 31896 30848 31932
rect 30884 31896 30924 31932
rect 30960 31898 31002 31932
rect 31036 31898 31076 31934
rect 30960 31896 31076 31898
rect 30818 31878 31076 31896
rect 31292 31932 31392 31968
rect 31292 31896 31324 31932
rect 31360 31896 31392 31932
rect 31292 31878 31392 31896
rect 30818 31804 31076 31822
rect 30818 31768 30848 31804
rect 30882 31768 30922 31804
rect 30956 31768 31002 31804
rect 31036 31768 31076 31804
rect 31292 31804 31392 31822
rect 31292 31768 31324 31804
rect 31360 31768 31392 31804
rect 30818 31732 31076 31768
rect 31292 31732 31392 31768
rect 30818 31662 31076 31696
rect 30818 31660 31002 31662
rect 30818 31624 30848 31660
rect 30884 31624 30924 31660
rect 30960 31626 31002 31660
rect 31036 31626 31076 31662
rect 30960 31624 31076 31626
rect 30818 31606 31076 31624
rect 31292 31660 31392 31696
rect 31292 31624 31324 31660
rect 31360 31624 31392 31660
rect 31292 31606 31392 31624
rect 30876 31474 31078 31492
rect 30876 31438 30918 31474
rect 30952 31438 31002 31474
rect 31036 31438 31078 31474
rect 30876 31402 31078 31438
rect 30876 31330 31078 31366
rect 30876 31294 30920 31330
rect 30956 31294 31002 31330
rect 31038 31294 31078 31330
rect 30876 31276 31078 31294
<< pdiff >>
rect 31610 33586 31868 33604
rect 31610 33550 31642 33586
rect 31678 33550 31714 33586
rect 31750 33550 31784 33586
rect 31820 33550 31868 33586
rect 31610 33514 31868 33550
rect 31610 33442 31868 33478
rect 31610 33406 31642 33442
rect 31678 33406 31712 33442
rect 31748 33406 31782 33442
rect 31818 33406 31868 33442
rect 31610 33388 31868 33406
rect 31610 33310 32186 33326
rect 31610 33308 31712 33310
rect 31610 33272 31642 33308
rect 31678 33274 31712 33308
rect 31748 33274 31782 33310
rect 31818 33274 31852 33310
rect 31888 33274 31922 33310
rect 31958 33274 31992 33310
rect 32028 33274 32062 33310
rect 32098 33274 32132 33310
rect 32168 33274 32186 33310
rect 31678 33272 32186 33274
rect 31610 33236 32186 33272
rect 31610 33164 32186 33200
rect 31610 33128 31642 33164
rect 31678 33128 31712 33164
rect 31748 33128 31782 33164
rect 31818 33128 31852 33164
rect 31888 33128 31922 33164
rect 31958 33128 31992 33164
rect 32028 33128 32062 33164
rect 32098 33128 32132 33164
rect 32168 33128 32186 33164
rect 31610 33110 32186 33128
rect 31610 32892 31710 32910
rect 31610 32856 31642 32892
rect 31678 32856 31710 32892
rect 31922 32894 32182 32912
rect 31922 32858 31964 32894
rect 31998 32858 32044 32894
rect 32078 32858 32118 32894
rect 32152 32858 32182 32894
rect 31610 32820 31710 32856
rect 31922 32822 32182 32858
rect 31610 32748 31710 32784
rect 31610 32712 31642 32748
rect 31678 32712 31710 32748
rect 31610 32694 31710 32712
rect 31922 32752 32182 32786
rect 31922 32716 31964 32752
rect 31998 32750 32182 32752
rect 31998 32716 32040 32750
rect 31922 32714 32040 32716
rect 32076 32714 32116 32750
rect 32152 32714 32182 32750
rect 31922 32696 32182 32714
rect 31610 32620 31710 32638
rect 31610 32584 31642 32620
rect 31678 32584 31710 32620
rect 31922 32622 32182 32640
rect 31922 32586 31964 32622
rect 31998 32586 32044 32622
rect 32078 32586 32118 32622
rect 32152 32586 32182 32622
rect 31610 32548 31710 32584
rect 31922 32550 32182 32586
rect 31610 32476 31710 32512
rect 31610 32440 31642 32476
rect 31678 32440 31710 32476
rect 31610 32422 31710 32440
rect 31922 32480 32182 32514
rect 31922 32444 31964 32480
rect 31998 32478 32182 32480
rect 31998 32444 32040 32478
rect 31922 32442 32040 32444
rect 32076 32442 32116 32478
rect 32152 32442 32182 32478
rect 31922 32424 32182 32442
rect 31610 32348 31710 32366
rect 31610 32312 31642 32348
rect 31678 32312 31710 32348
rect 31922 32350 32182 32368
rect 31922 32314 31964 32350
rect 31998 32314 32044 32350
rect 32078 32314 32118 32350
rect 32152 32314 32182 32350
rect 31610 32276 31710 32312
rect 31922 32278 32182 32314
rect 31610 32204 31710 32240
rect 31610 32168 31642 32204
rect 31678 32168 31710 32204
rect 31610 32150 31710 32168
rect 31922 32208 32182 32242
rect 31922 32172 31964 32208
rect 31998 32206 32182 32208
rect 31998 32172 32040 32206
rect 31922 32170 32040 32172
rect 32076 32170 32116 32206
rect 32152 32170 32182 32206
rect 31922 32152 32182 32170
rect 31608 32076 31708 32094
rect 31608 32040 31640 32076
rect 31676 32040 31708 32076
rect 31922 32078 32182 32096
rect 31922 32042 31964 32078
rect 31998 32042 32044 32078
rect 32078 32042 32118 32078
rect 32152 32042 32182 32078
rect 31608 32004 31708 32040
rect 31922 32006 32182 32042
rect 31608 31932 31708 31968
rect 31608 31896 31640 31932
rect 31676 31896 31708 31932
rect 31608 31878 31708 31896
rect 31922 31936 32182 31970
rect 31922 31900 31964 31936
rect 31998 31934 32182 31936
rect 31998 31900 32040 31934
rect 31922 31898 32040 31900
rect 32076 31898 32116 31934
rect 32152 31898 32182 31934
rect 31922 31880 32182 31898
rect 31608 31804 31708 31822
rect 31608 31768 31640 31804
rect 31676 31768 31708 31804
rect 31922 31806 32182 31824
rect 31922 31770 31964 31806
rect 31998 31770 32044 31806
rect 32078 31770 32118 31806
rect 32152 31770 32182 31806
rect 31608 31732 31708 31768
rect 31922 31734 32182 31770
rect 31608 31660 31708 31696
rect 31608 31624 31640 31660
rect 31676 31624 31708 31660
rect 31608 31606 31708 31624
rect 31922 31664 32182 31698
rect 31922 31628 31964 31664
rect 31998 31662 32182 31664
rect 31998 31628 32040 31662
rect 31922 31626 32040 31628
rect 32076 31626 32116 31662
rect 32152 31626 32182 31662
rect 31922 31608 32182 31626
rect 31922 31474 32124 31490
rect 31922 31472 32024 31474
rect 31922 31436 31954 31472
rect 31990 31438 32024 31472
rect 32060 31438 32124 31474
rect 31990 31436 32124 31438
rect 31922 31400 32124 31436
rect 31922 31328 32124 31364
rect 31922 31292 31964 31328
rect 32000 31292 32046 31328
rect 32082 31292 32124 31328
rect 31922 31274 32124 31292
<< ndiffc >>
rect 31326 33550 31362 33586
rect 31326 33406 31362 33442
rect 31132 33272 31166 33308
rect 31206 33272 31240 33308
rect 31274 33272 31308 33308
rect 31344 33272 31380 33308
rect 31132 33128 31166 33164
rect 31206 33128 31240 33164
rect 31274 33128 31308 33164
rect 31342 33128 31378 33164
rect 30848 32856 30882 32892
rect 30922 32856 30956 32892
rect 31002 32856 31036 32892
rect 31326 32856 31362 32892
rect 30848 32712 30884 32748
rect 30924 32712 30960 32748
rect 31002 32714 31036 32750
rect 31326 32712 31362 32748
rect 30848 32584 30882 32620
rect 30922 32584 30956 32620
rect 31002 32584 31036 32620
rect 31326 32584 31362 32620
rect 30848 32440 30884 32476
rect 30924 32440 30960 32476
rect 31002 32442 31036 32478
rect 31326 32440 31362 32476
rect 30848 32312 30882 32348
rect 30922 32312 30956 32348
rect 31002 32312 31036 32348
rect 31326 32312 31362 32348
rect 30848 32168 30884 32204
rect 30924 32168 30960 32204
rect 31002 32170 31036 32206
rect 31326 32168 31362 32204
rect 30848 32040 30882 32076
rect 30922 32040 30956 32076
rect 31002 32040 31036 32076
rect 31324 32040 31360 32076
rect 30848 31896 30884 31932
rect 30924 31896 30960 31932
rect 31002 31898 31036 31934
rect 31324 31896 31360 31932
rect 30848 31768 30882 31804
rect 30922 31768 30956 31804
rect 31002 31768 31036 31804
rect 31324 31768 31360 31804
rect 30848 31624 30884 31660
rect 30924 31624 30960 31660
rect 31002 31626 31036 31662
rect 31324 31624 31360 31660
rect 30918 31438 30952 31474
rect 31002 31438 31036 31474
rect 30920 31294 30956 31330
rect 31002 31294 31038 31330
<< pdiffc >>
rect 31642 33550 31678 33586
rect 31714 33550 31750 33586
rect 31784 33550 31820 33586
rect 31642 33406 31678 33442
rect 31712 33406 31748 33442
rect 31782 33406 31818 33442
rect 31642 33272 31678 33308
rect 31712 33274 31748 33310
rect 31782 33274 31818 33310
rect 31852 33274 31888 33310
rect 31922 33274 31958 33310
rect 31992 33274 32028 33310
rect 32062 33274 32098 33310
rect 32132 33274 32168 33310
rect 31642 33128 31678 33164
rect 31712 33128 31748 33164
rect 31782 33128 31818 33164
rect 31852 33128 31888 33164
rect 31922 33128 31958 33164
rect 31992 33128 32028 33164
rect 32062 33128 32098 33164
rect 32132 33128 32168 33164
rect 31642 32856 31678 32892
rect 31964 32858 31998 32894
rect 32044 32858 32078 32894
rect 32118 32858 32152 32894
rect 31642 32712 31678 32748
rect 31964 32716 31998 32752
rect 32040 32714 32076 32750
rect 32116 32714 32152 32750
rect 31642 32584 31678 32620
rect 31964 32586 31998 32622
rect 32044 32586 32078 32622
rect 32118 32586 32152 32622
rect 31642 32440 31678 32476
rect 31964 32444 31998 32480
rect 32040 32442 32076 32478
rect 32116 32442 32152 32478
rect 31642 32312 31678 32348
rect 31964 32314 31998 32350
rect 32044 32314 32078 32350
rect 32118 32314 32152 32350
rect 31642 32168 31678 32204
rect 31964 32172 31998 32208
rect 32040 32170 32076 32206
rect 32116 32170 32152 32206
rect 31640 32040 31676 32076
rect 31964 32042 31998 32078
rect 32044 32042 32078 32078
rect 32118 32042 32152 32078
rect 31640 31896 31676 31932
rect 31964 31900 31998 31936
rect 32040 31898 32076 31934
rect 32116 31898 32152 31934
rect 31640 31768 31676 31804
rect 31964 31770 31998 31806
rect 32044 31770 32078 31806
rect 32118 31770 32152 31806
rect 31640 31624 31676 31660
rect 31964 31628 31998 31664
rect 32040 31626 32076 31662
rect 32116 31626 32152 31662
rect 31954 31436 31990 31472
rect 32024 31438 32060 31474
rect 31964 31292 32000 31328
rect 32046 31292 32082 31328
<< psubdiff >>
rect 30678 33322 30714 33346
rect 30678 33262 30714 33286
rect 30678 33046 30714 33070
rect 30678 32986 30714 33010
rect 30678 32704 30714 32728
rect 30678 32644 30714 32668
rect 30678 32430 30714 32454
rect 30678 32370 30714 32394
rect 30678 32158 30714 32182
rect 30678 32098 30714 32122
rect 30678 31888 30714 31912
rect 30678 31828 30714 31852
rect 30678 31566 30714 31590
rect 30678 31506 30714 31530
<< nsubdiff >>
rect 32284 33308 32320 33332
rect 32284 33248 32320 33272
rect 32284 33050 32320 33074
rect 32284 32990 32320 33014
rect 32284 32742 32320 32766
rect 32284 32682 32320 32706
rect 32284 32472 32320 32496
rect 32284 32412 32320 32436
rect 32284 32214 32320 32238
rect 32284 32154 32320 32178
rect 32276 31938 32326 31972
rect 32276 31902 32286 31938
rect 32322 31902 32326 31938
rect 32276 31874 32326 31902
rect 32286 31586 32322 31610
rect 32286 31526 32322 31550
<< psubdiffcont >>
rect 30678 33286 30714 33322
rect 30678 33010 30714 33046
rect 30678 32668 30714 32704
rect 30678 32394 30714 32430
rect 30678 32122 30714 32158
rect 30678 31852 30714 31888
rect 30678 31530 30714 31566
<< nsubdiffcont >>
rect 32284 33272 32320 33308
rect 32284 33014 32320 33050
rect 32284 32706 32320 32742
rect 32284 32436 32320 32472
rect 32284 32178 32320 32214
rect 32286 31902 32322 31938
rect 32286 31550 32322 31586
<< poly >>
rect 31240 33478 31266 33514
rect 31396 33490 31610 33514
rect 31396 33478 31490 33490
rect 31474 33454 31490 33478
rect 31526 33478 31610 33490
rect 31868 33478 31894 33514
rect 31526 33454 31542 33478
rect 31474 33440 31542 33454
rect 31486 33430 31530 33440
rect 31082 33200 31108 33236
rect 31396 33212 31610 33236
rect 31396 33200 31490 33212
rect 31474 33176 31490 33200
rect 31526 33200 31610 33212
rect 32186 33200 32212 33236
rect 31526 33176 31542 33200
rect 31474 33162 31542 33176
rect 31486 33152 31530 33162
rect 31122 32856 31166 32866
rect 31110 32842 31178 32856
rect 31110 32820 31126 32842
rect 30792 32784 30818 32820
rect 31076 32806 31126 32820
rect 31162 32806 31178 32842
rect 31834 32858 31878 32868
rect 31822 32844 31890 32858
rect 31076 32784 31178 32806
rect 31258 32784 31294 32820
rect 31394 32796 31610 32820
rect 31394 32784 31490 32796
rect 31474 32760 31490 32784
rect 31526 32784 31610 32796
rect 31710 32784 31746 32820
rect 31822 32808 31838 32844
rect 31874 32822 31890 32844
rect 31874 32808 31922 32822
rect 31822 32786 31922 32808
rect 32182 32786 32208 32822
rect 31526 32760 31542 32784
rect 31474 32746 31542 32760
rect 31486 32736 31530 32746
rect 31122 32584 31166 32594
rect 31110 32570 31178 32584
rect 31110 32548 31126 32570
rect 30792 32512 30818 32548
rect 31076 32534 31126 32548
rect 31162 32534 31178 32570
rect 31834 32586 31878 32596
rect 31822 32572 31890 32586
rect 31076 32512 31178 32534
rect 31258 32512 31294 32548
rect 31394 32524 31610 32548
rect 31394 32512 31490 32524
rect 31474 32488 31490 32512
rect 31526 32512 31610 32524
rect 31710 32512 31746 32548
rect 31822 32536 31838 32572
rect 31874 32550 31890 32572
rect 31874 32536 31922 32550
rect 31822 32514 31922 32536
rect 32182 32514 32208 32550
rect 31526 32488 31542 32512
rect 31474 32474 31542 32488
rect 31486 32464 31530 32474
rect 31122 32312 31166 32322
rect 31110 32298 31178 32312
rect 31110 32276 31126 32298
rect 30792 32240 30818 32276
rect 31076 32262 31126 32276
rect 31162 32262 31178 32298
rect 31834 32314 31878 32324
rect 31822 32300 31890 32314
rect 31076 32240 31178 32262
rect 31258 32240 31294 32276
rect 31394 32252 31610 32276
rect 31394 32240 31490 32252
rect 31474 32216 31490 32240
rect 31526 32240 31610 32252
rect 31710 32240 31746 32276
rect 31822 32264 31838 32300
rect 31874 32278 31890 32300
rect 31874 32264 31922 32278
rect 31822 32242 31922 32264
rect 32182 32242 32208 32278
rect 31526 32216 31542 32240
rect 31474 32202 31542 32216
rect 31486 32192 31530 32202
rect 31122 32040 31166 32050
rect 31110 32026 31178 32040
rect 31110 32004 31126 32026
rect 30792 31968 30818 32004
rect 31076 31990 31126 32004
rect 31162 31990 31178 32026
rect 31834 32042 31878 32052
rect 31822 32028 31890 32042
rect 31076 31968 31178 31990
rect 31256 31968 31292 32004
rect 31392 31980 31608 32004
rect 31392 31968 31488 31980
rect 31472 31944 31488 31968
rect 31524 31968 31608 31980
rect 31708 31968 31744 32004
rect 31822 31992 31838 32028
rect 31874 32006 31890 32028
rect 31874 31992 31922 32006
rect 31822 31970 31922 31992
rect 32182 31970 32208 32006
rect 31524 31944 31540 31968
rect 31472 31930 31540 31944
rect 31484 31920 31528 31930
rect 31122 31768 31166 31778
rect 31110 31754 31178 31768
rect 31110 31732 31126 31754
rect 30792 31696 30818 31732
rect 31076 31718 31126 31732
rect 31162 31718 31178 31754
rect 31834 31770 31878 31780
rect 31822 31756 31890 31770
rect 31076 31696 31178 31718
rect 31256 31696 31292 31732
rect 31392 31708 31608 31732
rect 31392 31696 31488 31708
rect 31472 31672 31488 31696
rect 31524 31696 31608 31708
rect 31708 31696 31744 31732
rect 31822 31720 31838 31756
rect 31874 31734 31890 31756
rect 31874 31720 31922 31734
rect 31822 31698 31922 31720
rect 32182 31698 32208 31734
rect 31524 31672 31540 31696
rect 31472 31658 31540 31672
rect 31484 31648 31528 31658
rect 31122 31438 31166 31448
rect 31110 31424 31178 31438
rect 31834 31436 31878 31446
rect 31110 31402 31126 31424
rect 30850 31366 30876 31402
rect 31078 31388 31126 31402
rect 31162 31388 31178 31424
rect 31078 31366 31178 31388
rect 31822 31422 31890 31436
rect 31822 31386 31838 31422
rect 31874 31400 31890 31422
rect 31874 31386 31922 31400
rect 31822 31364 31922 31386
rect 32124 31364 32150 31400
<< polycont >>
rect 31490 33454 31526 33490
rect 31490 33176 31526 33212
rect 31126 32806 31162 32842
rect 31490 32760 31526 32796
rect 31838 32808 31874 32844
rect 31126 32534 31162 32570
rect 31490 32488 31526 32524
rect 31838 32536 31874 32572
rect 31126 32262 31162 32298
rect 31490 32216 31526 32252
rect 31838 32264 31874 32300
rect 31126 31990 31162 32026
rect 31488 31944 31524 31980
rect 31838 31992 31874 32028
rect 31126 31718 31162 31754
rect 31488 31672 31524 31708
rect 31838 31720 31874 31756
rect 31126 31388 31162 31424
rect 31838 31386 31874 31422
<< locali >>
rect 31310 33590 31394 33602
rect 31490 33590 31526 33630
rect 31610 33590 31860 33602
rect 31310 33586 31860 33590
rect 31310 33550 31326 33586
rect 31362 33550 31642 33586
rect 31678 33550 31714 33586
rect 31750 33550 31784 33586
rect 31820 33550 31860 33586
rect 31310 33546 31860 33550
rect 31310 33534 31394 33546
rect 31610 33534 31860 33546
rect 30656 33456 30734 33500
rect 31474 33490 31542 33500
rect 31306 33456 31378 33458
rect 30656 33444 31378 33456
rect 31474 33454 31490 33490
rect 31526 33454 31542 33490
rect 32262 33458 32336 33472
rect 31474 33446 31542 33454
rect 30656 33408 30678 33444
rect 30714 33442 31378 33444
rect 30714 33408 31326 33442
rect 30656 33406 31326 33408
rect 31362 33406 31378 33442
rect 30656 33394 31378 33406
rect 30656 33322 30734 33394
rect 31306 33390 31378 33394
rect 30656 33286 30678 33322
rect 30714 33286 30734 33322
rect 30656 33180 30734 33286
rect 31124 33312 31394 33324
rect 31490 33312 31526 33446
rect 31622 33442 32336 33458
rect 31622 33406 31642 33442
rect 31678 33406 31712 33442
rect 31748 33406 31782 33442
rect 31818 33406 32282 33442
rect 32318 33406 32336 33442
rect 31622 33390 32336 33406
rect 31610 33320 31692 33324
rect 31610 33312 32184 33320
rect 31124 33310 32184 33312
rect 31124 33308 31712 33310
rect 31124 33272 31132 33308
rect 31166 33272 31206 33308
rect 31240 33272 31274 33308
rect 31308 33272 31344 33308
rect 31380 33272 31642 33308
rect 31678 33274 31712 33308
rect 31748 33274 31782 33310
rect 31818 33274 31852 33310
rect 31888 33274 31922 33310
rect 31958 33274 31992 33310
rect 32028 33274 32062 33310
rect 32098 33274 32132 33310
rect 32168 33274 32184 33310
rect 31678 33272 32184 33274
rect 31124 33268 32184 33272
rect 31124 33258 31394 33268
rect 31132 33256 31394 33258
rect 31610 33256 32184 33268
rect 32262 33308 32336 33390
rect 32262 33272 32284 33308
rect 32320 33272 32336 33308
rect 31474 33212 31542 33222
rect 30656 33164 31392 33180
rect 31474 33176 31490 33212
rect 31526 33176 31542 33212
rect 32262 33182 32336 33272
rect 32164 33180 32336 33182
rect 31474 33168 31542 33176
rect 30656 33158 31132 33164
rect 30656 33122 30678 33158
rect 30714 33128 31132 33158
rect 31166 33128 31206 33164
rect 31240 33128 31274 33164
rect 31308 33128 31342 33164
rect 31378 33128 31392 33164
rect 30714 33122 31392 33128
rect 30656 33114 31392 33122
rect 30656 33112 31378 33114
rect 30656 33046 30734 33112
rect 30656 33010 30678 33046
rect 30714 33010 30734 33046
rect 30656 32906 30734 33010
rect 31490 32964 31526 33168
rect 31622 33166 32336 33180
rect 31622 33164 32282 33166
rect 31622 33128 31642 33164
rect 31678 33128 31712 33164
rect 31748 33128 31782 33164
rect 31818 33128 31852 33164
rect 31888 33128 31922 33164
rect 31958 33128 31992 33164
rect 32028 33128 32062 33164
rect 32098 33128 32132 33164
rect 32168 33130 32282 33164
rect 32318 33130 32336 33166
rect 32168 33128 32336 33130
rect 31622 33114 32336 33128
rect 31622 33112 32178 33114
rect 32262 33050 32336 33114
rect 32262 33014 32284 33050
rect 32320 33014 32336 33050
rect 30818 32906 31062 32908
rect 30656 32892 31062 32906
rect 30656 32890 30848 32892
rect 30656 32854 30678 32890
rect 30714 32856 30848 32890
rect 30882 32856 30922 32892
rect 30956 32856 31002 32892
rect 31036 32856 31062 32892
rect 30714 32854 31062 32856
rect 30656 32842 31062 32854
rect 31126 32850 31162 32884
rect 31310 32896 31394 32908
rect 31490 32896 31526 32922
rect 31610 32896 31692 32908
rect 31310 32892 31692 32896
rect 31310 32856 31326 32892
rect 31362 32856 31642 32892
rect 31678 32856 31692 32892
rect 31310 32852 31692 32856
rect 32262 32912 32336 33014
rect 32178 32910 32336 32912
rect 31838 32852 31874 32886
rect 31938 32906 32336 32910
rect 31938 32896 32338 32906
rect 31938 32894 32282 32896
rect 31938 32858 31964 32894
rect 31998 32858 32044 32894
rect 32078 32858 32118 32894
rect 32152 32860 32282 32894
rect 32318 32860 32338 32896
rect 32152 32858 32338 32860
rect 30656 32704 30734 32842
rect 30818 32840 31062 32842
rect 31110 32842 31178 32850
rect 31110 32806 31126 32842
rect 31162 32806 31178 32842
rect 31310 32840 31394 32852
rect 31610 32840 31692 32852
rect 31822 32844 31890 32852
rect 31822 32808 31838 32844
rect 31874 32808 31890 32844
rect 31938 32844 32338 32858
rect 31938 32842 32182 32844
rect 31110 32796 31178 32806
rect 31474 32796 31542 32806
rect 31822 32798 31890 32808
rect 30656 32668 30678 32704
rect 30714 32668 30734 32704
rect 30818 32754 31076 32766
rect 30818 32752 31078 32754
rect 31306 32752 31378 32764
rect 31474 32760 31490 32796
rect 31526 32760 31542 32796
rect 31474 32752 31542 32760
rect 31622 32754 31694 32764
rect 31924 32756 32182 32768
rect 31922 32754 32182 32756
rect 31622 32752 32182 32754
rect 30818 32750 31378 32752
rect 30818 32748 31002 32750
rect 30818 32712 30848 32748
rect 30884 32712 30924 32748
rect 30960 32714 31002 32748
rect 31036 32748 31378 32750
rect 31036 32714 31326 32748
rect 30960 32712 31326 32714
rect 31362 32712 31378 32748
rect 30818 32706 31378 32712
rect 30818 32696 31076 32706
rect 31306 32696 31378 32706
rect 30656 32634 30734 32668
rect 30818 32634 31062 32636
rect 30656 32620 31062 32634
rect 30656 32584 30848 32620
rect 30882 32584 30922 32620
rect 30956 32584 31002 32620
rect 31036 32584 31062 32620
rect 30656 32570 31062 32584
rect 31126 32578 31162 32612
rect 31310 32624 31394 32636
rect 31490 32624 31526 32752
rect 31622 32748 31964 32752
rect 31622 32712 31642 32748
rect 31678 32716 31964 32748
rect 31998 32750 32182 32752
rect 31998 32716 32040 32750
rect 31678 32714 32040 32716
rect 32076 32714 32116 32750
rect 32152 32714 32182 32750
rect 31678 32712 32182 32714
rect 31622 32708 32182 32712
rect 31622 32696 31694 32708
rect 31924 32698 32182 32708
rect 32262 32742 32338 32844
rect 32262 32706 32284 32742
rect 32320 32706 32338 32742
rect 31610 32624 31692 32636
rect 31310 32620 31692 32624
rect 31310 32584 31326 32620
rect 31362 32584 31642 32620
rect 31678 32584 31692 32620
rect 31310 32580 31692 32584
rect 32262 32640 32338 32706
rect 32180 32638 32338 32640
rect 31838 32580 31874 32614
rect 31938 32622 32338 32638
rect 31938 32586 31964 32622
rect 31998 32586 32044 32622
rect 32078 32586 32118 32622
rect 32152 32586 32284 32622
rect 32320 32586 32338 32622
rect 30656 32534 30678 32570
rect 30714 32534 30734 32570
rect 30818 32568 31062 32570
rect 31110 32570 31178 32578
rect 30656 32430 30734 32534
rect 31110 32534 31126 32570
rect 31162 32534 31178 32570
rect 31310 32568 31394 32580
rect 31610 32568 31692 32580
rect 31822 32572 31890 32580
rect 31822 32536 31838 32572
rect 31874 32536 31890 32572
rect 31938 32572 32338 32586
rect 31938 32570 32182 32572
rect 31110 32524 31178 32534
rect 31474 32524 31542 32534
rect 31822 32526 31890 32536
rect 30656 32394 30678 32430
rect 30714 32394 30734 32430
rect 30818 32482 31076 32494
rect 30818 32480 31078 32482
rect 31306 32480 31378 32492
rect 31474 32488 31490 32524
rect 31526 32488 31542 32524
rect 31474 32480 31542 32488
rect 31622 32482 31694 32492
rect 31924 32484 32182 32496
rect 31922 32482 32182 32484
rect 31622 32480 32182 32482
rect 30818 32478 31378 32480
rect 30818 32476 31002 32478
rect 30818 32440 30848 32476
rect 30884 32440 30924 32476
rect 30960 32442 31002 32476
rect 31036 32476 31378 32478
rect 31036 32442 31326 32476
rect 30960 32440 31326 32442
rect 31362 32440 31378 32476
rect 30818 32434 31378 32440
rect 30818 32424 31076 32434
rect 31306 32424 31378 32434
rect 30656 32364 30734 32394
rect 30656 32348 31062 32364
rect 30656 32312 30848 32348
rect 30882 32312 30922 32348
rect 30956 32312 31002 32348
rect 31036 32312 31062 32348
rect 30656 32300 31062 32312
rect 31126 32306 31162 32340
rect 31310 32352 31394 32364
rect 31490 32352 31526 32480
rect 31622 32476 31964 32480
rect 31622 32440 31642 32476
rect 31678 32444 31964 32476
rect 31998 32478 32182 32480
rect 31998 32444 32040 32478
rect 31678 32442 32040 32444
rect 32076 32442 32116 32478
rect 32152 32442 32182 32478
rect 31678 32440 32182 32442
rect 31622 32436 32182 32440
rect 31622 32424 31694 32436
rect 31924 32426 32182 32436
rect 32262 32472 32338 32572
rect 32262 32436 32284 32472
rect 32320 32436 32338 32472
rect 31610 32352 31692 32364
rect 31310 32348 31692 32352
rect 31310 32312 31326 32348
rect 31362 32312 31642 32348
rect 31678 32312 31692 32348
rect 31310 32308 31692 32312
rect 32262 32366 32338 32436
rect 31838 32308 31874 32342
rect 31938 32350 32338 32366
rect 31938 32314 31964 32350
rect 31998 32314 32044 32350
rect 32078 32314 32118 32350
rect 32152 32314 32286 32350
rect 32322 32314 32338 32350
rect 30656 32294 30734 32300
rect 30818 32296 31062 32300
rect 31110 32298 31178 32306
rect 30656 32258 30678 32294
rect 30714 32258 30734 32294
rect 30656 32158 30734 32258
rect 31110 32262 31126 32298
rect 31162 32262 31178 32298
rect 31310 32296 31394 32308
rect 31610 32296 31692 32308
rect 31822 32300 31890 32308
rect 31822 32264 31838 32300
rect 31874 32264 31890 32300
rect 31938 32298 32338 32314
rect 31110 32252 31178 32262
rect 31474 32252 31542 32262
rect 31822 32254 31890 32264
rect 30656 32122 30678 32158
rect 30714 32122 30734 32158
rect 30818 32210 31076 32222
rect 30818 32208 31078 32210
rect 31306 32208 31378 32220
rect 31474 32216 31490 32252
rect 31526 32216 31542 32252
rect 31474 32208 31542 32216
rect 31622 32210 31694 32220
rect 31924 32212 32182 32224
rect 31922 32210 32182 32212
rect 31622 32208 32182 32210
rect 30818 32206 31378 32208
rect 30818 32204 31002 32206
rect 30818 32168 30848 32204
rect 30884 32168 30924 32204
rect 30960 32170 31002 32204
rect 31036 32204 31378 32206
rect 31036 32170 31326 32204
rect 30960 32168 31326 32170
rect 31362 32168 31378 32204
rect 30818 32162 31378 32168
rect 30818 32152 31076 32162
rect 31306 32152 31378 32162
rect 31490 32160 31526 32208
rect 30656 32090 30734 32122
rect 31488 32132 31526 32160
rect 31622 32204 31964 32208
rect 31622 32168 31642 32204
rect 31678 32172 31964 32204
rect 31998 32206 32182 32208
rect 31998 32172 32040 32206
rect 31678 32170 32040 32172
rect 32076 32170 32116 32206
rect 32152 32170 32182 32206
rect 31678 32168 32182 32170
rect 31622 32164 32182 32168
rect 31622 32152 31694 32164
rect 31924 32154 32182 32164
rect 32262 32214 32338 32298
rect 32262 32178 32284 32214
rect 32320 32178 32338 32214
rect 30818 32090 31062 32092
rect 30656 32076 31062 32090
rect 30656 32040 30848 32076
rect 30882 32040 30922 32076
rect 30956 32040 31002 32076
rect 31036 32040 31062 32076
rect 30656 32026 31062 32040
rect 31126 32034 31162 32068
rect 31308 32080 31392 32092
rect 31488 32080 31524 32132
rect 31608 32080 31690 32092
rect 31308 32076 31690 32080
rect 31308 32040 31324 32076
rect 31360 32040 31640 32076
rect 31676 32040 31690 32076
rect 31308 32036 31690 32040
rect 32262 32094 32338 32178
rect 31838 32036 31874 32070
rect 31938 32080 32338 32094
rect 31938 32078 32286 32080
rect 31938 32042 31964 32078
rect 31998 32042 32044 32078
rect 32078 32042 32118 32078
rect 32152 32044 32286 32078
rect 32322 32044 32338 32080
rect 32152 32042 32338 32044
rect 30656 32022 30734 32026
rect 30818 32024 31062 32026
rect 31110 32026 31178 32034
rect 30656 31986 30678 32022
rect 30714 31986 30734 32022
rect 30656 31888 30734 31986
rect 31110 31990 31126 32026
rect 31162 31990 31178 32026
rect 31308 32024 31392 32036
rect 31608 32024 31690 32036
rect 31822 32028 31890 32036
rect 31822 31992 31838 32028
rect 31874 31992 31890 32028
rect 31938 32026 32338 32042
rect 31110 31980 31178 31990
rect 31472 31980 31540 31990
rect 31822 31982 31890 31992
rect 30656 31852 30678 31888
rect 30714 31852 30734 31888
rect 30818 31938 31076 31950
rect 30818 31936 31078 31938
rect 31304 31936 31376 31948
rect 31472 31944 31488 31980
rect 31524 31944 31540 31980
rect 31472 31936 31540 31944
rect 31620 31938 31692 31948
rect 31924 31940 32182 31952
rect 31922 31938 32182 31940
rect 31620 31936 32182 31938
rect 30818 31934 31376 31936
rect 30818 31932 31002 31934
rect 30818 31896 30848 31932
rect 30884 31896 30924 31932
rect 30960 31898 31002 31932
rect 31036 31932 31376 31934
rect 31036 31898 31324 31932
rect 30960 31896 31324 31898
rect 31360 31896 31376 31932
rect 30818 31890 31376 31896
rect 30818 31880 31076 31890
rect 31304 31880 31376 31890
rect 30656 31818 30734 31852
rect 30818 31818 31062 31820
rect 30656 31804 31062 31818
rect 30656 31768 30848 31804
rect 30882 31768 30922 31804
rect 30956 31768 31002 31804
rect 31036 31768 31062 31804
rect 30656 31754 31062 31768
rect 31126 31762 31162 31796
rect 31308 31808 31392 31820
rect 31488 31808 31524 31936
rect 31620 31932 31964 31936
rect 31620 31896 31640 31932
rect 31676 31900 31964 31932
rect 31998 31934 32182 31936
rect 31998 31900 32040 31934
rect 31676 31898 32040 31900
rect 32076 31898 32116 31934
rect 32152 31898 32182 31934
rect 31676 31896 32182 31898
rect 31620 31892 32182 31896
rect 31620 31880 31692 31892
rect 31924 31882 32182 31892
rect 32262 31938 32338 32026
rect 32262 31902 32286 31938
rect 32322 31902 32338 31938
rect 31608 31808 31690 31820
rect 31308 31804 31690 31808
rect 31308 31768 31324 31804
rect 31360 31768 31640 31804
rect 31676 31768 31690 31804
rect 31308 31764 31690 31768
rect 32262 31824 32338 31902
rect 32182 31822 32338 31824
rect 31838 31764 31874 31798
rect 31938 31808 32338 31822
rect 31938 31806 32286 31808
rect 31938 31770 31964 31806
rect 31998 31770 32044 31806
rect 32078 31770 32118 31806
rect 32152 31772 32286 31806
rect 32322 31772 32338 31808
rect 32152 31770 32338 31772
rect 30656 31710 30734 31754
rect 30818 31752 31062 31754
rect 31110 31754 31178 31762
rect 30656 31674 30678 31710
rect 30714 31674 30734 31710
rect 31110 31718 31126 31754
rect 31162 31718 31178 31754
rect 31308 31752 31392 31764
rect 31608 31752 31690 31764
rect 31822 31756 31890 31764
rect 31822 31720 31838 31756
rect 31874 31720 31890 31756
rect 31938 31756 32338 31770
rect 31938 31754 32182 31756
rect 32262 31754 32338 31756
rect 31110 31708 31178 31718
rect 31472 31708 31540 31718
rect 31822 31710 31890 31720
rect 30656 31566 30734 31674
rect 30818 31666 31076 31678
rect 30818 31664 31078 31666
rect 31304 31664 31376 31676
rect 31472 31672 31488 31708
rect 31524 31672 31540 31708
rect 31472 31664 31540 31672
rect 31620 31666 31692 31676
rect 31924 31668 32182 31680
rect 31922 31666 32182 31668
rect 31620 31664 32182 31666
rect 30818 31662 31376 31664
rect 30818 31660 31002 31662
rect 30818 31624 30848 31660
rect 30884 31624 30924 31660
rect 30960 31626 31002 31660
rect 31036 31660 31376 31662
rect 31036 31626 31324 31660
rect 30960 31624 31324 31626
rect 31360 31624 31376 31660
rect 30818 31618 31376 31624
rect 30818 31608 31076 31618
rect 31304 31608 31376 31618
rect 31488 31630 31524 31664
rect 31620 31660 31964 31664
rect 31620 31624 31640 31660
rect 31676 31628 31964 31660
rect 31998 31662 32182 31664
rect 31998 31628 32040 31662
rect 31676 31626 32040 31628
rect 32076 31626 32116 31662
rect 32152 31626 32182 31662
rect 31676 31624 32182 31626
rect 31620 31620 32182 31624
rect 31620 31608 31692 31620
rect 31924 31610 32182 31620
rect 30656 31530 30678 31566
rect 30714 31530 30734 31566
rect 30656 31484 30734 31530
rect 32264 31586 32338 31754
rect 32264 31550 32286 31586
rect 32322 31550 32338 31586
rect 30876 31484 31058 31490
rect 30656 31474 31058 31484
rect 30656 31472 30918 31474
rect 30656 31436 30678 31472
rect 30714 31438 30918 31472
rect 30952 31438 31002 31474
rect 31036 31438 31058 31474
rect 30714 31436 31058 31438
rect 30656 31430 31058 31436
rect 31126 31432 31162 31466
rect 32264 31484 32338 31550
rect 30656 31370 30734 31430
rect 30876 31422 31058 31430
rect 31110 31424 31178 31432
rect 31838 31430 31874 31464
rect 31934 31474 32338 31484
rect 31934 31472 32024 31474
rect 31934 31436 31954 31472
rect 31990 31438 32024 31472
rect 32060 31468 32338 31474
rect 32060 31438 32286 31468
rect 31990 31436 32286 31438
rect 31934 31432 32286 31436
rect 32322 31432 32338 31468
rect 31110 31388 31126 31424
rect 31162 31388 31178 31424
rect 31110 31378 31178 31388
rect 31822 31422 31890 31430
rect 31822 31386 31838 31422
rect 31874 31386 31890 31422
rect 31934 31420 32338 31432
rect 31822 31376 31890 31386
rect 30876 31336 31058 31348
rect 31828 31340 31878 31376
rect 31926 31340 32106 31344
rect 31828 31336 32106 31340
rect 30876 31330 32106 31336
rect 30876 31294 30920 31330
rect 30956 31294 31002 31330
rect 31038 31328 32106 31330
rect 31038 31294 31964 31328
rect 30876 31292 31964 31294
rect 32000 31292 32046 31328
rect 32082 31292 32106 31328
rect 30876 31284 32106 31292
rect 30876 31278 31058 31284
rect 31828 31282 32106 31284
rect 31922 31276 32106 31282
rect 32264 31186 32338 31420
rect 32264 30996 32336 31186
rect 32266 30830 32336 30996
rect 32266 30792 32282 30830
rect 32320 30792 32336 30830
rect 32266 30782 32336 30792
<< viali >>
rect 31490 33630 31526 33666
rect 30678 33408 30714 33444
rect 32282 33406 32318 33442
rect 30678 33122 30714 33158
rect 32282 33130 32318 33166
rect 31490 32922 31526 32964
rect 30678 32854 30714 32890
rect 31126 32884 31162 32922
rect 31838 32886 31874 32924
rect 32282 32860 32318 32896
rect 31126 32612 31162 32650
rect 31838 32614 31874 32652
rect 32284 32586 32320 32622
rect 30678 32534 30714 32570
rect 31126 32340 31162 32378
rect 31838 32342 31874 32380
rect 32286 32314 32322 32350
rect 30678 32258 30714 32294
rect 31126 32068 31162 32106
rect 31838 32070 31874 32108
rect 32286 32044 32322 32080
rect 30678 31986 30714 32022
rect 31126 31796 31162 31834
rect 31838 31798 31874 31836
rect 32286 31772 32322 31808
rect 30678 31674 30714 31710
rect 31488 31588 31524 31630
rect 30678 31436 30714 31472
rect 31126 31466 31162 31504
rect 31838 31464 31874 31502
rect 32286 31432 32322 31468
rect 32282 30792 32320 30830
<< metal1 >>
rect 31474 33820 31544 33900
rect 31470 33810 31548 33820
rect 31470 33754 31482 33810
rect 31538 33754 31548 33810
rect 31470 33734 31548 33754
rect 31478 33666 31536 33734
rect 30660 33582 30730 33662
rect 31478 33630 31490 33666
rect 31526 33630 31536 33666
rect 31478 33600 31536 33630
rect 30656 33572 30734 33582
rect 30656 33516 30668 33572
rect 30724 33516 30734 33572
rect 30656 33500 30734 33516
rect 30654 33496 30734 33500
rect 30654 33444 30736 33496
rect 30654 33408 30678 33444
rect 30714 33408 30736 33444
rect 30654 33158 30736 33408
rect 30654 33122 30678 33158
rect 30714 33122 30736 33158
rect 30654 32890 30736 33122
rect 32266 33442 32338 33470
rect 32266 33406 32282 33442
rect 32318 33406 32338 33442
rect 32266 33166 32338 33406
rect 32266 33130 32282 33166
rect 32318 33130 32338 33166
rect 31478 32964 31536 32976
rect 30654 32854 30678 32890
rect 30714 32854 30736 32890
rect 30654 32570 30736 32854
rect 30654 32534 30678 32570
rect 30714 32534 30736 32570
rect 30654 32294 30736 32534
rect 30654 32258 30678 32294
rect 30714 32258 30736 32294
rect 30654 32022 30736 32258
rect 30654 31986 30678 32022
rect 30714 31986 30736 32022
rect 30654 31710 30736 31986
rect 30654 31674 30678 31710
rect 30714 31674 30736 31710
rect 30654 31472 30736 31674
rect 30654 31436 30678 31472
rect 30714 31436 30736 31472
rect 30654 31368 30736 31436
rect 31116 32922 31174 32936
rect 31116 32884 31126 32922
rect 31162 32884 31174 32922
rect 31116 32650 31174 32884
rect 31116 32612 31126 32650
rect 31162 32612 31174 32650
rect 31116 32378 31174 32612
rect 31116 32340 31126 32378
rect 31162 32340 31174 32378
rect 31116 32106 31174 32340
rect 31116 32068 31126 32106
rect 31162 32068 31174 32106
rect 31116 31834 31174 32068
rect 31116 31796 31126 31834
rect 31162 31796 31174 31834
rect 31116 31504 31174 31796
rect 31116 31466 31126 31504
rect 31162 31466 31174 31504
rect 31116 31438 31174 31466
rect 31478 32922 31490 32964
rect 31526 32922 31536 32964
rect 31478 31630 31536 32922
rect 31478 31588 31488 31630
rect 31524 31588 31536 31630
rect 31116 31366 31226 31438
rect 31478 31088 31536 31588
rect 31826 32924 31884 32938
rect 31826 32886 31838 32924
rect 31874 32886 31884 32924
rect 31826 32652 31884 32886
rect 31826 32614 31838 32652
rect 31874 32614 31884 32652
rect 31826 32380 31884 32614
rect 31826 32342 31838 32380
rect 31874 32342 31884 32380
rect 31826 32108 31884 32342
rect 31826 32070 31838 32108
rect 31874 32070 31884 32108
rect 31826 31836 31884 32070
rect 31826 31798 31838 31836
rect 31874 31798 31884 31836
rect 31826 31502 31884 31798
rect 32266 32896 32338 33130
rect 32266 32860 32282 32896
rect 32318 32860 32338 32896
rect 32266 32622 32338 32860
rect 32266 32586 32284 32622
rect 32320 32586 32338 32622
rect 32266 32350 32338 32586
rect 32266 32314 32286 32350
rect 32322 32314 32338 32350
rect 32266 32080 32338 32314
rect 32266 32044 32286 32080
rect 32322 32044 32338 32080
rect 32266 31808 32338 32044
rect 32266 31772 32286 31808
rect 32322 31772 32338 31808
rect 32266 31748 32338 31772
rect 31826 31464 31838 31502
rect 31874 31464 31884 31502
rect 31826 31364 31884 31464
rect 32264 31468 32338 31748
rect 32264 31432 32286 31468
rect 32322 31432 32338 31468
rect 32264 31368 32338 31432
rect 32208 31088 32462 31090
rect 31478 31084 32602 31088
rect 31478 31076 32682 31084
rect 31478 31020 32536 31076
rect 32592 31020 32682 31076
rect 31478 31014 32682 31020
rect 32516 31010 32602 31014
rect 32268 30830 32334 30846
rect 32268 30792 32282 30830
rect 32320 30792 32334 30830
rect 32268 30784 32334 30792
rect 32272 30736 32330 30784
rect 32260 30716 32338 30736
rect 32260 30660 32270 30716
rect 32326 30660 32338 30716
rect 32260 30650 32338 30660
rect 32264 30570 32334 30650
<< via1 >>
rect 31482 33754 31538 33810
rect 30668 33516 30724 33572
rect 32536 31020 32592 31076
rect 32270 30660 32326 30716
<< metal2 >>
rect 31474 33820 31544 33900
rect 31470 33810 31548 33820
rect 31470 33754 31482 33810
rect 31538 33754 31548 33810
rect 31470 33734 31548 33754
rect 30660 33582 30730 33662
rect 30656 33572 30734 33582
rect 30656 33516 30668 33572
rect 30724 33516 30734 33572
rect 30656 33496 30734 33516
rect 32516 31084 32602 31088
rect 32516 31076 32682 31084
rect 32516 31020 32536 31076
rect 32592 31020 32682 31076
rect 32516 31014 32682 31020
rect 32516 31010 32602 31014
rect 32260 30716 32338 30736
rect 32260 30660 32270 30716
rect 32326 30660 32338 30716
rect 32260 30650 32338 30660
rect 32264 30570 32334 30650
<< via2 >>
rect 31482 33754 31538 33810
rect 30668 33516 30724 33572
rect 32536 31020 32592 31076
rect 32270 30660 32326 30716
<< metal3 >>
rect -5555 48669 -5275 48743
rect -5347 34018 -5277 48669
rect 40745 45713 40815 48711
rect -5346 33853 -5277 34018
rect 31474 45650 40815 45713
rect 31474 45643 39644 45650
rect -5346 33783 30730 33853
rect 31474 33820 31544 45643
rect 30660 33582 30730 33783
rect 31470 33810 31548 33820
rect 31470 33754 31482 33810
rect 31538 33754 31548 33810
rect 31470 33734 31548 33754
rect 30656 33572 30734 33582
rect 30656 33516 30668 33572
rect 30724 33516 30734 33572
rect 30656 33496 30734 33516
rect 32516 31084 32602 31088
rect 32516 31076 52417 31084
rect 32516 31020 32536 31076
rect 32592 31020 52417 31076
rect 32516 31014 52417 31020
rect 32516 31010 32602 31014
rect 32260 30716 32338 30736
rect 32260 30660 32270 30716
rect 32326 30660 32338 30716
rect 32260 30650 32338 30660
rect 32264 30585 32334 30650
rect 32264 -11876 32335 30585
rect 52347 26995 52417 31014
rect 52347 26925 54401 26995
rect 32264 -11947 54145 -11876
<< end >>
